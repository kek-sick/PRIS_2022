En man i orange hatt stirrar på något.
En Boston Terrier kör på lummigt grönt gräs framför ett vitt staket.
En tjej i karateuniform som bryter en pinne med en framspark.
Fem personer med vinterjackor och hjälmar står i snön, med snöskotrar i bakgrunden.
Folk håller på att laga taket på ett hus.
En man i ljusa kläder fotograferar en grupp män som bär mörka kostymer och hattar som står runt en kvinna klädd i en axellös klänning.
En grupp människor som står framför en igloo.
En pojke i röd uniform försöker undvika att komma ut på hemmaplan, medan fångvaktaren i den blå uniformen försöker fånga honom.
En kille jobbar på en byggnad.
En man i väst sitter i en stol och håller i tidningar.
En mor och hennes unga sång njuter av en vacker dag utanför.
Män som spelar volleyboll, med en spelare som saknar bollen men händerna fortfarande i luften.
En kvinna som håller en skål mat i ett kök.
Man sitter med verktyg vid ett bord i sitt hem.
Tre personer sitter i en grotta.
En flicka i jeansklänning går längs en höjd balansstråle.
En blondin som håller hand med en kille i sanden.
En kvinna i grå tröja och svart keps står i kö i en affär.
Personen i randig skjorta är bergsklättring.
Två män låtsas vara stadgar medan kvinnor ser på.
Folk står utanför en byggnad.
En tonåring spelar trumpet på planen på en match.
En kvinna gör en somersault på en studsmatta på stranden.
En man står vid en grupp videospel i en bar.
En kvinna använder en övning medan en annan man tar en bild.
En kvinna i rosa tröja och ett förkläde, som rengör ett bord med en svamp.
En man som hugger grenar av träd.
Grupp av asiatiska pojkar väntar på kött att laga mat över grillen.
Kvinnor, som bär traditionella kläder, återverkar sitt eget liv.
En man håller ner en annan mans huvud och förbereder sig för att slå honom i ansiktet.
Sex personer rider mountainbikes genom en djungelmiljö.
2 blonda tjejer sitter på en avsats i ett trångt torg.
Ett barn plaskar i vattnet
Tre personer sitter vid ett picknickbord utanför en byggnad målad som en fackjacka.
Tre pojkar står på en pir i sina baddräkter.
En anställd ger en kvinna en väska medan hon surfar genom fisk på is på en gatumarknad.
En vacker kvinna spelar harpsichord.
Utanför en byggnad tittar en uniformerad säkerhetsvakt på kameran bakom ett staket.
Den unga damen tittar på pizzan.
En skjortlös man i shorts fiskar medan han står på några klippor.
En flicka med flytväst flyter i vatten.
En man i uniform och en man i blå skjorta står framför en lastbil.
Folk sitter inne i ett tåg.
Ett barn svänger med fötterna uppe i luften i en skog.
En man i röd skjorta går in på en anläggning.
Två män som bär badbyxor hoppar upp i luften på en måttligt befolkad strand.
Ett litet barn lagar mat med en annan person.
En fader-figur och två barn utanför deras hem gör gårdsarbete som att använda en hoe på gräset och plantera ett träd.
En man som lagar mat på spisen.
En man i jeans på stranden som leker med en röd boll.
Folk går längs trottoaren bredvid en rad butiker.
En wakeboarder utför en flip samtidigt bogseras i hög hastighet.
En stor grupp människor fyller en gata.
En man på en tagglinje som går ner i vattnet.
En kvinna i jeans går förbi en buss med en annons som skildrar en kvinna som kikar över sina solglasögon.
En man i rosa skjorta sitter i gräset och en boll är i luften.
En bil parkerad vid stranden.
Två män klädda i svart i en stad
Mannen i gula byxor höjer armarna.
Två män som bär hattar och använder käppar går nära en vattenförekomst under solnedgången.
Ett hejarklacksteam som gör en rutin på stolar.
En pojke spelar schack med en vuxen som visas utanför skärmen medan en flicka tittar på.
En massa människor ute för lite kul i den allmänna parken.
En man sitter på en bänk och håller sin hund och tittar på vattnet.
En pojke och hans yngre bror leker tillsammans på lekplatsen.
En kvinna i blått ser i en svart läderväska medan hon sitter på en bänk under en solig eftermiddag medan människor och limousiner passerade bakom henne.
Den bruna hunden står på sandstranden.
En kvinna sitter med en korg tyg, omgiven av tyg.
En man grillar ute på sin bakgård.
En kvinna sjunger i en klubb med en gitarrist bakom sig.
Gitarrspelaren uppträder på en nattklubbsröd gitarr.
Ett barn som sitter på en gräsmatta och tittar upp mot kameran
Två damer och tre män som tittar på havet.
En kvinnlig artist med violin spelar på en gata medan en kvinna med en blå gitarr tittar på.
En ung flicka som simmar i en pool
Flera barn är utomhus och gör sig redo att leka dragkamp.
Tre tonåringar i en tunnelbana leker runt.
En brun hund går i gräset med tungan hängande ut.
Folk som sitter i gräset utanför en byggnad och tar en paus.
Tröjlös kille stirrar iväg på avstånd medan tre kvinnor går förbi en publik som sitter utanför ett café.
Två unga pojkar som sätter frukt på cykeln.
En man i svart t-shirt, keps och jeans spelar trummor på en upp och ner gul pail.
En ung kvinnlig konstnär målar en bild av en kvinna på en vägg.
Två kvinnliga medlemmar i laget USA utför ett hopp high-fem omgiven av två andra kvinnliga medlemmar.
En man som rör om i en kruka med vätska i det här köket.
Pojken vaknar på sjön.
En man jobbar på ett korvstånd.
En stor grupp människor i olika åldrar och kön sitter utanför tillsammans.
En blondhårig kvinna häller drinkar på en bar.
Ett litet barn bär en blå och vit t-shirt glatt håller en gul plast alligator.
En kvinna med rosa hår klädd i svart pratar med en man.
Mannen i japansk matlagningsdräkt förbereder en måltid för två personer.
En flicka hoppar över floden, från sten till sten.
En manlig arbetare med sin verktygslåda knäböjer bredvid två kvinnor.
En äldre man öppnar sina armar vida och ser förbryllad ut.
Ett barn i en vit karate outfit övar ett drag
Tre män i samma färgade västar är utomhus.
En kvinna tar en bild av ett barn som bär en rosa hatt medan en man bär henne.
En grupp mest asiatiska barn som sitter på bås i blå stolar.
En ung pojke i en fotbollsuniform som gråter i sina handflator.
En lycklig kvinna förbereder en förfriskning på ett kafé.
En byggnadsarbetare kör tung utrustning på en arbetsplats.
En kvinna springer efter att ha gjort en träff i kvinnors softball, fångaren stiger till hennes fötter.
En man i arbetsuniform som skickar ett verktyg till en annan person.
En grupp människor klättrar i kallt väder.
En bergsklättrare som är på väg nerför ett berg med en blå hjälm på.
En man som står på en rund staty.
Ett barn som sitter vid ett restaurangbord och håller en pappersmask mot ansiktet.
En brun hund vadar in i en sjö för att hämta en pinne.
En mor lär sina två unga pojkar att fiska utanför en stenig kust i mycket blått vatten.
Ett litet barn går bredvid röda banderoller.
En flicka sitter på en dekorerad cykel med en yngre pojke medan en annan flicka tar en bild.
En svart hund hämtar en boll i vatten.
En man i vita byxor och en blå skjorta sparkar en gul boxningssäck.
Två indianer deltar i en ceremoni.
En pojke med en skadad näsa och skrivande på händerna står i en videouthyrningsbutik.
Två siluettmänniskor paddlar en kanot på havet under solnedgången.
Människor står på en fullsatt tunnelbana, och plattformen utanför syns genom fönstret.
Människan skalvägg med eld i handen
Två bruna hundar springer genom snön.
På scen foto av små band uppträda för teater publik.
En bebis i juldräkt tittar på kameran.
En man sitter bredvid en datormonitor.
Den här damen har hört ett roligt skämt och skratta.
Människor inne i en byggnad, en tar ett foto.
Fyra vita hundar med mynningar hoppar över en röd vägg.
Kvinnan med den blå skjortan håller i ett barn.
Två personer sitter och fiskar på randiga strandstolar i en vattenförekomst.
En gammal kvinna som jobbar i en vävstol och tillverkar tyg.
En pojke som står i förgrunden och ser ut över andra människor i en domstol.
En man i en blå rock som tar en ung pojkes axel.
Tre bruna hundar hoppar upp mot kvinnan i blått.
En pojke hänger ut ur en förbipasserande taxi taxi fönster
En man i grå skjorta hoppar över toppen av en sanddyn i öknen.
Ett barn som bär gul skjorta hoppar upp och ner.
En arbetare i gul jacka lyfts upp högt för att arbeta på en byggnad.
En man i Brasilien höll ett informellt tal med unga vuxna.
En massa öl drar flikar i en bar med julbelysning i taket.
En man är på väg nerför en klippa över havet.
En svart man går till sin lastbil i snön.
En rävterrier hoppar efter en boll.
En kvinnlig polis i en mössa och marin uniform ler medan han bär solglasögon utanför en butik.
En familj går en promenad i en park.
En man i grön hård hatt och gul skyddsväst rynkar.
Barn med rosa strängar på huvudet dansar omgiven av konfetti, ballonger.
En hund med en snobbnäsa luktar för något på en flodbank.
En man förbereder sin lokala monter för dagarnas affärer.
En man i röd skjorta ska precis äta en taco.
En ung dam i vitt som håller i ett tennisracket
En pojke som bär en röd skjorta gräver i sanden med en gul spade.
En enskild bär rosenjacka plats sysslolös på en trä bänk.
En man som bär vit skjorta tittar ut genom ett fönster av en metallkonstruktion.
En kvinna håller i en liten vit staty.
Sex skjortlösa barn leker i naturligt vatten och plaskar runt.
Två personer cyklar genom en bergig region.
En flicka hoppar rep på en trottoar nära ett parkeringsgarage.
En man i orange skjorta och hjälm.
En liten pojke leker med plastblock, bilar och djur med en vuxen som tittar noga.
En liten flicka som öppnar en julklapp.
Kvinnan i blått har en kamera framför två andra kvinnor.
En liten flicka försöker ta en tupplur på den bekväma soffan.
En brun och svart hund som springer på en stig i skogen.
Två hundar leker vid ett träd.
En marin som går i svart rock och byxor på trappan när kameran fokuserar på hunden
Två män klädda i grönt lagar mat på en restaurang.
En man klädd i svart läder och en cowboyhatt går runt på en renässansfestival.
En hund springer ut med en gul leksak.
En hund som bär ett täcke springer i snön.
En familj leker på stranden med sin hund.
En kvinna och ett barn omfamnar medan barnet smakar vad de har gjort.
Två män och en dam står utanför.
En grupp män som använder stockar för att skjuta upp en båt ur vattnet.
En man dricker ur ett vinglas medan han läser tidningen.
En man klädd i svart och spelar piano.
En ung pojke med blå jersey och gula shorts spelar fotboll.
En man står på en stenstruktur med armarna ut som en fågel.
En hund dricker vatten ute på gräset.
Två kvinnor med tanklock tittar på kameran.
En man sitter i en frisörstol och gör sig redo för rakning.
Ett ungt barn som bär gröna stövlar och leker i en lerpöl
En man som använder en motorsåg för att hugga virke.
En man som satt vid ett picknickbord med en bricka och delvis drack öl framför sig.
Pojken med svart skjorta och blå jeans håller i ett rött basebollträ.
En mörkhårig skäggig man i glasögon och en Hawaiisk skjorta sitter på gräset.
Hundar springer på en hundkapplöpningsbana.
En lätt tekniker man med stamtatueringar som riktar en spotlight över en balkong.
Två tyska sheperder snyftar på varandra.
Detta är en grupp människor som står runt någon form av händelse.
En brun och vit hund som hämtar en leksak.
En man med vitt hår som spelar dragspel mitt i vissa byggnader.
En kvinna med brunt hår som sitter på en bänk utanför ett café.
En man bredvid en cykel spelar panflöjt.
Två barn balanserar på en stock och håller i ett rep.
En man som kör motorcykel utför ett trick på ett spår.
En ung kvinna med en lila duk som döljer hennes ansikte slappnar av på ett trädäck.
Kvinnan i den bruna skjortan sitter på en ljusröd bänk.
En hund går på en stock över en liten flod.
En ung man i vit t-shirt och gröna och svarta shorts står på en stubbe.
Alla människor är täckta av paraplyer.
En man annonserar med en stor skylt fastbunden på sin cykel.
En man kastar en stock i en vattenväg medan två hundar tittar.
De äldste spelar instrument under ett tält vid vattnet.
En utsikt över en fullsatt stadsgata.
En ung blond kvinna håller i ett vitt rep en solig dag.
Två personer i blå skjortor är ute med en bullhorn.
En svart hund dyker upp i en pool.
En cowboy rider på baksidan av en bronco i en tävling.
En järnvägsarbetare utför underhåll på järnvägsspår.
En arbetare i orange väst använder en spade.
Två byggnadsarbetare har en diskussion på arbetsplatsen.
Tre män går uppför kullen.
En asiatisk kvinna i en blommig bröllopsklänning poserar på en bro nära sina tärnor.
En ung man sjunger sin gitarr i köket.
Tre pojkar leker med svamp och hinkar med vatten.
Tre byggnadsarbetare lagar trottoaren.
Folk kyler ner sig i skogen bredvid kanoter.
En körgrupp samlas i en kyrka.
En grupp unga tonåringar hoppar på natten och gör roliga poser för kameran.
Två killar paddlar kajak, en orange en blå, nerför en bäck.
Två arbetare spred cement på en tegelbyggnad.
En dam med röd tröja och jeans sitter med händerna på vänster knä
Två artister sätter på en hånfull kamp för en publik som tittar uppmärksamt.
En GI slappnar av och väntar på en flygplats.
En man i gul rock tar hand om en brand, en pojke i en parka tittar.
En man och en pojke på en stenig strand.
En kvinna på en båt som heter "El Corazon" sänker svarta vikter i vattnet.
En pojke som sitter på och ser ut från ett mikroskop.
En ung barfota flicka i rosa klänning hoppar ut.
Många sitter runt ett tält utanför.
En ungdom med en svart skjorta som säger "Asien Pacific 2007" spelar en trumma när man sitter.
En man som säljer föremål nära vägkanten till det stora berget Canyon.
Flickan i gult skrattar åt flickan i orange medan hon blir bevakad av flickan i blått.
En hund hoppar över ett hinder utanför.
Hund med svart krage rullar i smuts och torkade blad
Två bruna hundar spelar på ett tufft sätt.
En man med mustasch och skägg håller i en stekpanna som har lågor som stiger från den.
En man, som bär revolutionerande menskläder, ringer en klocka.
En man i svart skjorta som fiskar på en stenig strand.
Två hundar är förbryllande varandra nos till nos.
Två män stannar för att prata på trottoaren när en bil passerar förbi.
En kinesisk man som sitter och väntar på kunder.
Parkerade bilar med en skolbuss bakom sig.
Två kvinnor med liknande skjortor går till vänster.
Ett litet barn bär en orange livväst som håller en åra paddling en blå kajak i en vattenförekomst.
Folk går på en stig i en trädfylld park.
Tre unga vuxna pratar i en skara människor, kvinnan ser upprörd ut.
Kvinna och barn utanför dörren till deras natursköna hem.
En svart man och hans två vita vänner håller ihop sina huvuden.
En tjej med kamouflagebyxor sitter ovanpå en Hummer.
En ljusbrun hund är på väg.
En pojke poserar med en stor grön insekt på näsan.
En skallig man demoniserar hur högt hans bruna och svarta hund kan hoppa.
En folksamling på en upptagen dagtid gata.
En greyhoundhund i gult och svart springer på banan.
En man som bär sandaler sitter på trottoaren nära några väskor.
En man och en kvinna sitter på basen av stängsel och har ett samtal.
Ett barn tittar på kaffemaskiner i en affär.
En man som dricker ur en gul kopp runt folk vid en hektisk händelse
En pojke lutar sig mot en bil med blommor på huven.
En kvinna i blommig klänning pratar med barn framför en skåpbil.
En man på sin bröllopsdag.
En ung kvinna med svart skjorta och jeans svepande.
Kvinna med hatt på att klättra på en klippa nära en stor vattenförekomst.
En stor svart pudel som springer på gräset med en leksak i munnen.
En shortspojke som gör ett skateboardtrick.
En liten pojke klädd i röda byxor står på gatan.
En kvinna sms på sin telefon, omgiven av paraplyer.
Åtta män spelar instrument på scenen, med en gitarrist framhävd i ljus.
En man i orange overall och matchande hård hatt hjälper till med en blå slang
En man och två flickor visar upp en fisk medan de håller fiskestolpar framför en vattenförekomst.
Man i röd skjorta tittar på hund på en agility kurs.
En pojke som bär röda och vita badbyxor dyker baklänges i en vacker pool.
En asiatisk kvinna som tar tillbaka håret.
En äldre kvinna och ett litet barn i en rosa skjorta som leker med flerfärgade block.
En liten svart hund hoppar över portarna
En brunhårig man i grön skjorta spelar trumpet utomhus.
En man pratar i telefon med fötterna uppe.
En grupp barn sitter på en blå matta medan de äter ur skålar.
En svart pojke sitter i sanden.
En liten hund tittar på två stora hundar som spelar hårt på ett fält.
Folk som sitter i en cirkel utanför en stor byggnad.
En hund hoppar för att fånga en softball medan en annan ser på.
Ett blond barn som svänger på en gunga.
En man och två kvinnor har en diskussion om vitt vin
En asiatisk man lagar mat utomhus.
En brun hund som ska fånga en grön frisbee.
Fans hejar när bandet spelar en låt.
En ung pojke står bredvid en sandskulptur av en pyramid.
Tre små barn går genom en gräsbevuxen trädgård.
En man lägger kilo på ett konstverk på en vagn.
En man på en cykel rider på ett berg.
En pojke med blå och gula regnstövlar springer på smuts.
En kvinna i orange jacka sitter på en bänk.
En man som gör ett trick på skateboard
En man i kampsportsuniform i luften.
En kvinna som säljer fruktpåsar på trottoaren.
Två fotbollslag är på planen.
Ett barn i en blå skjorta som hoppar från en bänk.
En målvakt i ett gult fält skyddar målet.
En grupp ungdomar skjuter i en mexikansk miljö.
En ung man åker skateboard från ett rosa räcke.
En ung pojke hoppar från en våningssäng på en mindre säng.
Två personer som bär udda alienliknande dräkter, en blå och en lila, står på en väg.
Man springer med en blå skjorta med ett nummer tejpat på.
En asiatisk fabriksarbetare poserar för kameran.
En man som verkar springa i ett maraton ger oss 2 tummar upp.
Basketspelare skjuter för ett mål under ett spel.
En fotbollsspelare i orange uniform ler och håller i fotbollen.
Två nedförsbacke skateboardåkare runt en kurva medan andra tittar.
Ett lag i vitt och guld vid sidan av en fotbollsplan.
En liten flicka knuffar sin skoter genom ett gräsrött trädkantat fält.
Grupp av asiatiska barn klädda i vita skjortor och hattar som uppträder med en publik som tittar på.
Fotgängare som går nerför gatan tittar på ett barn i en kartong.
En brun hund springer nerför sandstranden.
Två män i arméuniform står bredvid en kvinna.
Dali Lama under en mottagning där deltagarna har tagit med sig nejlikor, parasoller och böneflaggor.
En cyklist hoppar ett hinder.
Ett par sitter i vita gräsmatta stolar ler mot kameran.
Unga barn är på en liten tågresa.
En surfare i en blå baddräkt rider på vågorna.
Pojken hoppar på sin fotbollsspelare bror.
Två unga män på motsatta fotbollslag tävlar för att få bollen på en fotbollsplan.
Människor går på en asfalterad sluttning omgiven av kinesiska försäljare.
En ung pojke med vita byxor hoppar från soffan.
En pojke i orange skjorta häller legos ur en väska.
Kvinnan bär bruna sandaler och blå jeans, i en vit skjorta, håller ett barn under ett högt träd.
Tre människor ler och håller politiska tecken.
En polis står bredvid en bil på en stadsgata.
Två män i hatt.
En pojke i luften som försöker sparka en fotboll
En ung pojke med blå mössa har huvudet nere.
En rödhårig man med dreadlocks sitter och spelar och akustisk gitarr.
En man som äter en smörgås med sin dotter i knät.
Ett afrikanskt amerikanskt barn håller upp något som de i bilden är stolta över.
En kvinna leder en skara människor med en högtalare.
Utrustade åskådare ser på när en uniformerad polis håller ett tal och en man i kostym håller en skål med frukt.
En publik är närvarande på en bar.
En flicka i vitt och en flicka i grönt går förbi en blå biltvätt station.
En man använder elektronisk utrustning.
En person som surfar genom en kraschande våg i havet.
En officer inspekterar något.
En brud och brudgummen kysser under brudens slöja.
Riotpolisen står i bakgrunden medan en ung man med en röd halsduk som täcker hans ansikte går.
En svart och vit hund hoppar över ett brant valv i en tävling
En kvinna som bär tröja läser en bok i sitt hem.
Flera tonåringar tittar över ett räcke i ett mörkt rum.
Mannen i den vita t-shirten börjar klättra upp för en sten.
En tonårspojke stretchar i köket och man kan se en del av hans mage.
Människor håller olika typer av trumpinnar ovanför olika typer av trummor.
Tre jordbrukare skördar ris på ett risfält.
Två kvinnor och en man tittar på en bok.
Tre barns ben visas när de står nära en enda röra av fåniga snören.
En kock poserar för en kamera medan han lagar mat.
Många människor på en gata protesterar mot användningen av kol i kraftverk.
Tonåringen hoppar på kullen med sin cykel.
En liten flicka som springer på stranden.
Vit anka som flaxar sina vingar i vattnet.
Två män verkar samtala medan de står framför en lastbilsrygg och bakom ett metallföremål, medan fyra personer står runt dem.
En kvinna i rosa kjol håller i ett barn.
En hockeyspelare i en gul jersey vaktar målet.
En man går förbi en stor skylt som säger E.S.E. Electronics.
Tre pojkar med gröna skjortor och solbrända byxor poserar högst upp på en rutschkana.
En man dansar med en hund mellan benen.
Den vita hunden springer i det grunda vattnet.
Oregons slagverkare marscherar med bandet.
En grupp barn leker tillsammans på en inhägnad gård som en vuxen klocka.
En grupp kvinnor spelar musikinstrument tillsammans.
En liten flicka i en lila rutig klänning ligger på golvet och gråter.
En man med grått hår rakar skägget.
Två svarta hundar, en svart valp och en vit hund i snön.
En man i Miamis basketuniform som hoppar för att göra ett skott.
En kvinna sitter utanför sitt hus med en blå dörr och njuter av luften.
Ungar sitter på en man i banandräkt.
En grå och vit hund hoppar över stående vatten i sanden.
En folkmassa samlades runt en park vattenfontän i regnet.
Flera äldre män, några i traditionell huvudbonad samlas i ett gathörn.
En ung Lassie-hund är i snön.
Fotbollsspelaren som bär guldtröjan blockerar bollen från motståndarlagets spelare.
En kvinna i svart skjorta stickar med lila garn.
Fyra honor av asiatisk härkomst bär gyllene klänningar medan de utför punktbalett.
En person spelar ett unikt instrument.
En tjej som bär svarta sportkläder med nummer 1102 på sin tröja springer över lite gräs.
Ett barn längdskidor bär nummer "93".
En äldre gentleman och en ung flicka börjar arbeta på ett pussel tillsammans.
Ett filmteam filmar en ung afrikansk pojke i gul skjorta.
En gatubelysning upplyst bro med en cyklist och några bilar.
En man rider en tjur i en bullpen.
En pojke hoppar för att slå en tennisboll med sitt racket
Barn klättrar på en vägg som två andra tittar på.
Folk som går omkring på ett universitetsområde med palmer i bakgrunden.
Lilla flicka sparkar svart föremål på karate klass.
Två män som försöker lyfta sig upp från vattnet till en gångväg av däck.
Två män breakdancing, med en publik tittar på.
En professionellt klädd kvinna som står på ett podium och diskuterar något viktigt.
En kvinna ligger på en soffa och skrattar.
Ett jordgolv sopas av en vit och en svart kvinna.
En hjort hoppar över ett stängsel.
Tre hundar leker med varandra ute på fältet.
Två små barn ligger på sand.
En leende ung pojke leker i löven bland ankorna.
Dessa fyra personer står utomhus, med 3 hundar.
När man besöker Mayaruinerna pekar en guide i riktning mot fler attraktioner.
Tjejen som bär radio-t-shirt har öppen mun
En stamgrupp som fyller vattenkannor i öknen.
En man som står på en stadsgata.
En flock fåglar flyger iväg med mat i sina näbbar.
Två män rider genom åkermarken när de styr sin muledrivna trailer.
Två personer står på toppen av ett berg.
En ung flicka som roar sig när hon gör en snöängel.
Tre killar som ler mot kameran och visar upp sina muskler.
En person skriver på en krittavla i ett tomt klassrum.
En man i svart skjorta som sitter vid ett bord med en öppen Apple laptop framför sig.
Fyra personer slappnar av på en gräsbevuxen kulle med utsikt över en stenig dalgång.
En pojke med skateboard om han hoppar i luften längs några järnvägsspår.
Det finns en man i orange skjorta som spelar tennis.
Hunden med den röda kragen bär tänderna på hunden med den blå kragen.
Pojken är ute och njuter av en sommardag.
En arbetare i orange arbetsdräkt knäböjer och inspekterar en maskin.
Män i cowboyhattar står på en rodeo.
Det finns två hundar i snön och en har något i munnen.
En anställd tar en paus från arbetet för att ta en drink
En beige hund springer bakom en vit hund som håller en gul leksak.
Hockeyspelare i vit uniform med pinne
En man i vit skjorta med guldklocka som leker med ett kretskort.
En svart häst sticker huvudet genom ett stängsel och försöker nå gräset.
En crackhead låtsas hålla händerna varma men han röker faktiskt crack.
Två killar och en tjej som ler.
Ett barn lutar sig över en display som består av blå och gul plast, medan en vuxen tittar på.
En svartvit hund går för en tillplattad boll på snön.
En ung flicka som står bredvid en gul katt på en köksbänk.
De två barnen leker på lekplatsen.
En tennisspelare i en grön randig skjorta håller handen mot munnen.
En pojke i röd kostym leker i vattnet.
Ett barn som bär röd rock och mössa håller i en stor snöbit.
Två officerare med orangea jackor står utanför ett vitt tält med åskådare.
Två personer står bredvid ett träd på marken.
Två män sitter och pratar nära en stenbyggnad.
Ett brunettbarn med glasögon som håller ett blont barn i röd tröja och gula stövlar.
En svart och vit hund leker med en vit boll.
Två personer kysser varandra på en trottoar framför en limousin medan folk går förbi.
En kvinna spelar volleyboll.
Två stora hundar slåss på ett jordfält.
En brun hund hoppar över ett hinder.
En man i randig skjorta röker en cigarett på gatan
En liten flicka håller en liten pojke i knät.
En man som försöker rida en mycket galen tjur på en vacker lördag eftermiddag.
Barn slåss för att vinna en dragkamp.
En cyklist lutar en mountainbike runt en krök på en grusbana.
Två personer och en koppel ko på ett hem.
Den unge pojken lär sig cykla med sin pappa.
Pojke i röd skjorta och svarta shorts sopar uppfart.
En afrikansk familj står framför några provisoriska hus.
En man som spelar ett instrument bredvid ett träd.
Två kvinnor håller händerna över ett bord och ler mot kameran.
En flämtande brun hund som går på gräset.
En baseballspelare i en svart skjorta märkte just en spelare i en vit skjorta.
En kvinna håller en stor check på Kids Food Basket.
De två hundarna, en med en tennisboll i munnen, springer genom högt gräs.
Två vuxna och två barn sitter på en parkbänk.
En kvinna på ett gräsfält blåser på en maskros.
En man säljer potatis till en grupp människor.
En grupp människor på en gata samlas för att lyssna på ett dragspel.
En man sitter på en bänk lista till sin iPod
En gammal man på en tunnelbana som bär tunga kläder läser en tidning.
En äldre man i glasögon tillagar kött.
En man som utför ett trick på en cykel genom att stå på pedalerna medan cykeln är upprätt.
En man är på stranden och gör en sandskulptur.
Flera människor i en park äter vid ett picknickbord
Två kvinnor är fastspända vid ett träd i någon form av byggnadsarbete.
En cowboy i en rodeo som försöker slå klockan åtta.
En hund hoppar genom ett brinnande hinder.
En överviktig kvinna med långt svart hår i en rosa skjorta med namnbricka applicerar läppstift.
En man som fixar en liten flickas cykel.
Två flickor i puffiga kjolar dansar framför några musiker på gatan.
Den gula hunden bär en pinne med vatten.
En tjej i en tröja blockerar solstrålarna.
En rockkonsert äger rum.
Tre kvinnor i ljusa färger och huvudbonader håller kärlekskort.
En brun hund gräver i jorden.
Ung pojke i vit randig skjorta och pannband med tennisracket.
Två hundar springer iväg från kameran i skogen.
En flicka leker i fontänen påklädd.
Tre unga sumobrottare står och lyssnar på en kungörare
Två hanvandrare inspekterar en stock vid sidan av en skogsstig.
Tre spelare tar ett lag motståndare till marken.
Två pojkar går över en gata medan de sparkar en röd fotboll.
En man som håller upp en annan med ryggen.
Vit hund på bergssidan vänder sig mot något utanför scenen, himlen i bakgrunden.
En pojke som åker skateboard på en skateboardramp
En långhårig, manlig musiker spelar på ett piano.
Tre idrottare håller buketter står på seger podiet.
Två kala drag queens i röda klänningar
En ung pojke hänger på ett klädställ.
En liten flicka som bär rosa håller i en bar.
En man i grönt hoppar servermotorcyklar på sin egen motorcykel.
En kvinna som leker med två unga pojkar i en park
Fyra personer spelar fotboll på en strand.
Två tonårsflickor kramas, en bär cykelhjälm, med cyklister i bakgrunden.
Två medelstora hundar springer över snön.
En kvinna står på ett grönt fält och håller en vit hund och pekar på en brun hund.
Ett bord fullt av bilder i ramar, på en utomhusmarknad.
Två personer sitter vid ett bord utanför mot en vägg och gör ansikten.
Två killar med piercing i bröstvårtan ler.
Ett barn ligger på en beige matta och skrattar.
En man och kvinna är inlåsta armar som sitter ner och är uppklädda.
Två kvinnor brottas med lera i en barnpool.
En kille i vit skjorta går med en drink i handen.
Två personer är silhuetterade mot en sjö som reflekterar en målad himmel.
Flera personer sitter vid ett bord i formella kläder.
Två flickor (en klädd i blått och en klädd i rosa) tävlar varandra på rullskridskor.
De fyra människorna sitter på en hög med stenar.
En grupp människor gör tricks på motorcyklar.
Cyklist i racing redskap rider genom skogsområdet.
En man i grön skjorta går på stranden och bär sina gympaskor.
Flera män står runt en antik racerbil
Två män jobbar under huven på en vit racerbil.
Barn hoppar ner i en pool.
En man på kanten av en mur som håller på att ramla av.
En kvinna i randig klädsel på en cykel.
En flicka klädd i svart poserar för kameran.
Man i shorts står vid vattnet.
Fyra svarta män sitter på trappan till en kyrka.
En kran fungerar bland högar av spillror.
En gymnast klädd i rött och vitt är mitt-twirl på en ojämn bar.
En äldre dam i en grön tröja väljer grönsaker.
Två män tillverkar föremål i en verkstad med verktyg.
En lärare i vitt och en liten flicka i gul klänning som leker med byggsten.
Ett litet barn som sover i sängen med en öppen bok på bröstet.
En kvinna som äter i gräset en vacker dag.
En man går nerför en kullerstensgata bredvid byggnader målade solbränna med röda takrännor.
En kvinna som bär hatt och bakar bröd.
En ensam kvinna använder en stor primitiv murbruk och mortel för att krossa växtmaterial när hon står i ett stubbfält.
En man i karate uppträder inför två domare.
En man i formell klädsel spelar piano på trottoaren på en stadsgata.
En äldre man som sitter i en stol och äter lite snacks.
En kvinna i vit skjorta jobbar bakom disken på ett café.
En man med arbetskläder står på baksidan av en lastbil.
Två barn tittar på hästar genom ett litet staket.
Ett fönster med någon typ av design målad på den.
En kvinna som bär en ljusrosa ytterrock gör ett ansikte till en kvinna som bär en lila ytterrock medan hon står utanför en vitaminshoppa.
En cowboy slår ihop armen med ett bandage.
En man i gul skjorta och en man i mörkblå skjorta som pratar.
Tre asiatiska barn sitter på en soffa med gobelänger hängande i bakgrunden.
En tjej i röd skjorta hoppar upp för att träffa en tennisboll.
En man som poserar kameran med grön kran.
En man klinker flaskor med en annan person medan han ler på en restaurang.
En man lastar en låda lastbil med massor av bakade kringlor.
En man i svart jacka spelar gitarr offentligt.
En dansgrupp uppträder i en parad i Kina.
En man står på en klippa med utsikt över en vattensamling.
Polisen tittar på kvinnans utgång från bussen.
Två medelålders poliser vakar över en parkeringsplats på natten.
Två män i blå skjortor tittar på en fotbollsmatch.
En grupp män i blå uniformer står tillsammans.
En ung dam som gör yoga på stranden.
En stor skara människor står runt i en park och några spelar instrument.
En man med ballonghatt gör ballongdjur.
En man grillar kött på en grillgrop utomhus.
Två män säljer frukt på en fruktmarknad.
Brunettkvinna i en vit bikini som häller en drink i en mans kopp.
Pojke i solglasögon springer bakom en mässa.
En handskehänt hand håller vad som verkar vara en överdimensionerad nagel mot en stock.
En man i rutig skjorta visar upp en svart uppsättning handskar.
Två män i vita plaststolar sitter i en dörröppning.
En ung flicka i röd klänning bär en svart cowboyhatt.
Man i röd och vit fotboll uniform står på fältet gränslinjer med gul och blå fotboll.
Folk hoppar över en bergsspricka på ett rep.
Folk ser på som deltagare i ett maratonpass.
Människor på bärbara datorer framför pf ett stort fönster.
En diskjockey som är upptagen på jobbet när ljuset lyser på honom.
En man som bär handskar bär majs genom ett fält.
Ett foto är taget av en spegelreflektion av ett café.
En muslimsk kvinna som håller ballonger vid en islamisk händelse
En kvinna sitter i en bur i området med en katt och två kaniner.
En kvinna som sitter mot en tegelvägg inuti en byggnad.
Tre unga kvinnor möter varandra medan de sitter på röda plyschstolar.
En kvinna i blå skjorta som går i en by.
Sex barn som sitter på ett steg med anteckningsblock och kritor.
En brun hund som leker med en pinne på stranden.
Två hundar biter lekfullt en tredje hund, som har tungan stickande ut.
Ett barn är på en motorcykel och ler.
6 personer samlas runt för att äta en stor middag.
Jultomten fotograferas på ett evenemang.
Militärfamiljer marscherar genom New York en regnig dag.
En kvinna i blå hjälm och röda byxor som kör motorcykel.
Flera män bär kampsport uniformer medan de utför några drag i unisont.
En ung dam och man klädda i krigare kostym svinga pinnar med en grupp människor i bakgrunden.
En man i uniform går på en gata med två bilar och ett träd.
Ung kvinna klättrar rock ansikte
En äldre man i en ljusblå rock arbetar på en bil vid vägkanten.
Folk som tittar över flera färgade pappersbitar utspridda på ett bord.
En man sjunger och spelar gitarr i en mikrofon.
Två män sitter på en restaurang.
Två kvinnor i shorts springer nerför en strand längs vattnet.
Byggarbetare som har en diskussion vid spåren.
En utsikt över en gågata med en man i svart förkläde och en vit keps i mitten av bilden.
En grupp människor spelar på ett objekt.
En liten flicka i blå kläder klättrar på metallräcken på gatan.
En grupp män sitter och pratar bakom några gröna frukter.
En kille med gula kläder som står bakom en mikrofon under ett tält.
En brun hund med en lila frisbee i munnen.
Det ser ut som om en man som utövar sin kampsport rör sig nära ett lerigt vatten.
En kvinna med en drink och en kvinna med en mobiltelefon.
Ett barn i en röd rock viftar en hand i luften medan det ligger i snö bredvid en röd plastsläde.
En kvinna som sitter bredvid sin handväska och tittar på hundar i parken.
Tre män står på en scen, en bär clownmakeup och håller en gitarr.
En kvinna bearbetar växtvätska i en stamby
Kvinnan i den röda klänningen dansar med mannen i kostym.
Två små hundar följer en större hund med en tennisboll
En man med buskigt skägg och keps sitter på en parkbänk.
En afrikansk stam står i sin trädgård med skogen i bakgrunden.
En ung flicka försöker borsta en get.
Asiater sitter på en restaurang med gula stolar.
En liten flicka äter en kaka medan hon sitter i en barnstol och bär en haklapp.
En gråhårig man som bär svarta handskar flyttar gräsmattan.
En kvinna läser en bok medan hon sitter i en rad röda stolar.
Ett barn klappar medan det rider på en kvinnas axlar.
En familj går på trottoaren genom snön medan en man sitter på sidan med sin pappersmugg.
En katt sitter ovanpå en skylt.
En man i rosa skjorta och svart jacka med hörlurar på.
En ung man som ska kasta en fotboll.
En kille och en flicka som går längs en spiralväg.
En kvinna med rosa hår böjd ner på trottoaren håller för rosa hundar.
En man i kostym som håller en dryck i en kopp går längs trottoaren, bredvid en stadsbuss.
Man hoppar med en rockformation i bakgrunden.
En person i en röd jacka med svarta byxor som håller regnbågsband.
En kvinna lägger armen på en person som sitter i rullstol.
En man i ett vitt förkläde lagar något med ägg på en kastrull utanför för en kvinna i en solbränd jacka.
En kvinna med mobil och headset väntar på en korsning.
En grupp män går nerför en gata.
En väg bredvid en intressant plats med massor av pelare.
En grupp personer i svart står på en brygga i närheten en lång byggnad.
En man som bär några lådor öl.
En medelålders man sitter ner och spelar dragspel.
Tjej med grönt armband, hårband och örhängen står utanför.
En ung flicka i rosa skjorta är på en strand som springer mot havet.
En skateboardåkare i svart t-shirt och jeansåkning kastade staden.
En man i en jacka fotograferar en stor byggnad.
Folk vid sidan av en fotbollsmatch.
På det här fotot finns en familj på fyra personer som rusar över en livlig gata i staden.
En grupp människor går nerför gatan i solen.
En gata nära ett stoppljus med flera personer inklusive en man som bär en brun rock och solglasögon med handen mot ansiktet.
Vissa växter växer nära fönstret.
Denna spelare med den blå hjälmen var på slagträ och just avslutat svänger på bollen under ett lag baseball spel.
Kvinnan i guldrocken skyndar sig att fånga tunnelbanan.
En del människor sitter på bänkar under rader av träd framför en byggnad.
En man i kostym sitter vid en busshållplats.
En afrikansk amerikansk man omgiven av tomma vältade vita hinkar och mörkfärgade lådor uttrycker sig genom ett meddelande som är handskrivet på kartong.
En ung brunettkvinna som äter och dricker något.
En man i kostym och hatt spelar gitarr på gatan.
En kvinna i röd väst som jobbar på en dator.
Folk står runt rökelsen och viftar röken i ansiktet.
En man som använder badrumsspegeln för att knyta slipsen.
Musik spelas av flera individer medan en glad publik sitter och lyssnar.
Två unga män som rider på en mycket liten hästdragen vagn full av potatis.
En kvinna i klänning som går längs gatan förbi en byggarbetsplats.
En expedit i en närbutik frågar en kund som köper alkohol för sin ålder och identifiering.
En man med solglasögon kör en byggbil och släpper ut grus på marken.
En bebis som leker med sina leksaker och tittar på en svart och vit katt.
En tonårsflicka bär gitarr i skogen.
En man med ryggsäck går nerför gatan.
Två män har ett samtal framför en souvenirbutik i Rom.
En svart kvinna håller något i munnen.
En grupp människor sitter utomhus runt ett litet, kort bord.
En man som cyklar uppför rampen.
En kvinna som bär en svart tanktopp och ett korshalsband stirrar ut i fjärran nära solnedgången.
Tre unga flickor går tillsammans längs trottoaren.
En kvinna med långt hår är på en examensceremoni.
En man skateboardar på en väg medan en annan man tittar på från trottoaren.
En man i svart läderrock står framför en skylt.
En man och en kvinna som sjunger en sång tillsammans utanför.
En ung flicka med lockigt blont hår och bär en vit topp ligger i gräset, håller en blomma stjälk.
En ung dams fotbollslag med gröna uniformer utför en stretching motion.
En kvinna spelar ut en dramatisk scen offentligt bakom gult varningsband.
En man hukar sig medan han gör sysslor, när duvor vandrar i bakgrunden.
En grupp män som står på ett fält av svarta bollar.
En hektisk dag för medborgarna vid en lokal stadsdomstol.
En man med en cigarett i munnen som fixar en tallrik mat.
Två grupper simmare vadar ut.
Människor sitter på en bänk i en stad torg med slumpmässiga föremål inklusive en lampa och en klädskapare form stående i närheten.
Arbetarna omger ett hål med en hink.
En skjortlös man i svarta shorts står på den klippiga stranden till en stor vattenförekomst.
En vakt håller utkik medan han är i tjänst.
Folk spelar pool, en är en man som bär en blå skjorta och de andra är kvinnor men deras huvuden är inte inom kameran skott.
Folk står framför en skulptur omgiven av vatten.
En kvinna ser på som en man med vikta armar talar.
Medelålders man i vita shorts och flip-flops tittar upp på vägen
Två män klädda i mörk orange beläggningar och sandaler står nära en stor reflekterande skulptur.
Två personer tillbringar bra tid i sin båt.
En man och en kvinna står på gatan i staden.
Brandmän kommer från en tunnelbanestation.
Fyra män, av vilka tre bär bönemössor, sitter på en blå och olivgrön mönstrad matta.
Detta är en stor grupp människor som sitter utanför på bänkar.
En man i röd skjorta går förbi en turkos och vit rutig matinrättning som heter "32 De Neude".
Läkare som utför någon typ av operation.
En äldre man med en cigarett i munnen och en bollmössa inspekterar sin kamera.
Liten orkester som spelar med öppet violinfodral framför
En man med röd kostym dansar med en dam.
Två personer tittar på på natten vid lamporna i en stad.
Två motocross cyklister bär full skyddsutrustning, med en i luften efter ett hopp och den andra tittar ner på sin motorcykel.
Flera män klädda i orange samlas för en utomhus social händelse.
Två unga flickor springer på en trottoar utanför en tegelbyggnad med banderoller på.
Två enskilda klättrar upp för ett brant berg.
Ett barn ligger på marken bredvid en barnvagn.
En hund som tigger till en man och en kvinna.
Många människor på marknaden tittar på olika saker.
Två unga män spelar elgitarrer på scenen.
En tatuerad man häller öl ur en flaska i en ung mans mun.
Två personer står utanför och spränger leksaker och sopcontainrar.
Fyra personer cyklar på en cykelväg nära en livlig gata.
En kvinna i rosa skjorta och glasögon.
En kvinna i röd skjorta som lyfter armen till den förbipasserande folkmassan nedanför.
En pojke i vita shorts hoppar ner i en sjö eller flod.
En liten flicka tittar genom ett teleskop på stranden.
Flera byggnadsarbetare med orange skyddsvästar gräver ner i marken.
En person i en huva står framför en rasande byggnad.
Byggarbetare som picketar mot PM Construction Services.
En man som rider på en häst med några andra män som gör samma sak bakom sig.
En afroamerikansk man som gick nerför gatan.
Två nunnor poserar för en bild.
En kvinna med neonhörlurar skriver i en anteckningsbok.
En kvinna i grönmönstrad skjorta pratar på en mobiltelefon.
Ett litet afrikanskt barn bär ett yngre barn på ryggen.
En grupp människor sitter i stolar.
En person i en bandanna står på gatan framför sina saker.
En orientalisk person i röd skjorta och svarta byxor hukar sig över en handväska på betong.
En svart hund och en brun hund med boll.
En man med svart väst som håller ett modellflygplan
En man i ett fält med ett flygplan i sikte.
En man i kostym och slips och en kvinna med bagage förenar sig med andra i väntan på Londons tunnelbana.
Ett barn går längs trottoaren med några amerikanska flaggor.
En svart hund springer på grönt gräs med en leksak i munnen.
En orientalisk resenär väntar på sin tur vid valutaväxlingen.
En hund vänder sig mot gräset för att få fram en flygande boll.
En grupp elever sitter och lyssnar på talaren.
Folk kör scooters nerför gatan på natten.
En stor grå havsdäck och en kille på cykeln.
En man i orange skjorta och en blond pojke rider med andra människor på en "Pullman" fordon.
En ung man och kvinnor nära en stor metallskulptur
En båt med röda, vita och blå segel som dockar vid en brygga.
En man i svart hatt som fotograferar på en livlig gata.
En man står på en livlig gata och tittar med huvudet lutat uppåt.
En svart kvinna har en liten flicka i gul klänning på axlarna.
En grupp människor på gatan sätter upp instrument.
En fallen smutscyklist får hjälp av en annan.
Tre personer går uppför en bergsstig, medan en kvinna tittar på sin kamera.
Flera asiatiska män bär svarta kläder på någon form av station.
En kvinna i röd kjol går på gatan med graffiti i bakgrunden.
En rytmisk gymnast i en blå och rosa outfit utför en band rutin.
Folk svalkar i en fontän, en kvinna i vit klänning sitter på kanten och tittar på.
En man som sitter på en bänk under ett stort träd.
Tre män i röda och vita randiga skjortor, vita byxor och svarta hattar håller flaggor.
Folk beundrar ett konstverk.
Upptaget Asiatiskt köpcentrum med papperslyktor och shoppare.
Dessa människor klättrar uppför trappan för att gå till berget
Ett litet barn i blå kläder tittar bort på några träd i fjärran.
Folk tittar på barnleksaker i en affär.
En man med hatt spelar trummor på gatan.
En pojke står med tre flickor.
En leende man som bär ryggsäck håller upp nävarna framför en pojke i glasögon.
Fyra män är utanför och tittar ner över den gröna bron de är på.
En kvinna sover på en handduk framför folk som njuter av det blå vattnet.
En vuxen australiensisk herde följer efter en körande australiensisk herdevalp.
Fall shoppare och bistro mat älskare fångas i ebb och flöde av staden.
Den afroamerikanska mannen protesterar mot olagligt sex.
En polis är på en cykel och väntar på att ljuset ska bytas.
En grupp män sitter runt ett bord.
Högklassiga affärsmän inklusive äldre män har drinkar i parken.
Kvinna pratar med vän medan promenadhund ute på en solig dag.
En ung man i grå och svart skjorta och ett vitt pannband
Två personer kör motorcykel tillsammans med många andra förare.
Två kvinnor i militäruniform står med andra soldater i formation.
Tre flickor ler för en bild.
Damen med svarta fälgade glasögon och en gul tröja jacka ser förvirrad ut när hon sitter på solbränna täckt bänk.
En rödhårig ung man dricker ur en vattenfontän formad som en kvinna.
Två män och en kvinna går på en gata.
En medelålders man med rött hår och glasögon som håller ett spädbarn.
En ung pojke i röd hatt rider på en häst.
Två pojkar leker på trottoaren.
En liten flicka i svart baddräkt som håller en spade på en strand.
Gubben med hatt och kappa som sover uppe på en soffa.
Två pojkar tittar upp mot himlen och viftar med sina armar och de är klädda i kläder för att hålla dem varma.
Ett ungt par sitter på trottoaren och slappnar av tillsammans.
En ung man med skjorta och slips hukar sig ner och ger fredstecken.
Tre personer sitter vid ett bord utanför Bar Gelati Tabacchi.
En pojke i svart skjorta och röda armband hängande upp och ner medan andra människor tittar på.
En man som går framför en färgglad väggmålning.
En ung man som går med en annan ung man blickar tillbaka på tre flickor de just passerade
En man som putsar en palm inne i ett uteplats-liknande café'.
Fem personer gick uppför en trappa ledd av en kvinna i rosa skjorta och brun kjol.
En grupp människor på en marknad för frukt utomhus
Två pojkar äter sin McDonalds-lunch i en uteservering omgiven av många andra människor.
En kvinna som bär en jeansjacka går längs en trottoar
En man som kör ett fyrahjuligt fordon med fyra passagerare som rider fram och en man som sitter i sidled på baksidan.
En man i en tölpskjorta läser en tidning.
En pojke i barnvagn bär en grön skjorta och håller i en bok.
Två barn sitter sida vid sida medan de äter en godbit.
Folk cyklar på gatan, och de har alla hjälmar på sig.
Alla människor cyklar.
En man som sitter på en plattform med hjul dras av en håla.
En man på en cykel trampar genom en valvväg.
En färgglad ung man med synliga hudskador sitter och röker en cigarett.
Två män i kostym under paraply och framför graffiti.
En gammal mager man som bär den smutsiga vita skjortan och rider på en cykel på gatan
På hästryggen försöker en man repa en ung tjur.
En cowboy försöker lasso en kalv medan han rider en häst.
Två cykelister med hjälmar på rider förbi några tomma fält.
En man lutar sig över och drar upp något ur en påse.
En man i en bil åker förbi för att bevittna parkområdet.
En person med tatueringar tittar på ett foto på en digitalkamera, eller mobiltelefon.
En man i svart skjorta och jeans står på trottoaren och tittar på kameran.
En pojke och flicka står tillsammans på trottoaren när de tittar på ett föremål.
Flera personer i blå skrubb och en i kjol och svart blus.
En kvinna och en hund sitter på en vit bänk nära en strand.
Två kvinnor går i smuts utanför en stor byggnad.
En grupp män och ett barn i vita skjortor står på vägen.
En kvinna klädd i svart och bär en svart väska på trottoaren
Grupp av män som sitter runt ett bord och har ett samtal.
En väggmålning på sidan av en byggnad.
En asiatisk man som bär handskar arbetar på ett matstånd.
Kvinnan sitter vid ett bord medan hon arbetar på sin bärbara dator.
En person tittar på datorn på ett skrivbord med en telefon och en låda.
En man sitter i en stol och tittar på folk som går förbi.
Två människor som bär hattar står på ett fält och vårdar en gröda.
Vissa hoppar över en hög bar i Barcelona.
En man klädd i stövlar och en cowboyhatt sitter ovanpå en häst som hoppar medan åskådare sitter i läktaren.
Två unga flickor sitter på gatan och äter majs.
Tre barn i fotboll uniformer i två olika lag spelar fotboll på en fotbollsplan, medan en annan spelare och en vuxen står i bakgrunden.
Ett litet barn med ett smutsigt ansikte som hålls av en gammal kvinna.
En man med glasögon tittar på kameran medan en annan man i en blå skjorta tittar uppmärksamt på något.
Två personer som sitter under ett träd och plockar en grön grönsak.
En ung pojke med blå hatt tittar genom ett teleskop medan en annan pojke tittar.
3 män lagar mat i ett litet kök.
En ung flicka i grå snödräkt som åker skidor på ett snöigt berg.
En grupp bykvinnor samlades i dans
En man och en kvinna sorterar genom tvätt med latexhandskar på.
En ung flicka som sitter på en trästol.
Två arbetare svetsade galler på ett stängsel nära en livlig förortsgata.
En långhårig ung man som åker skateboard på rälsen en molnig dag.
På en utomhusmarknad skyfflar två män snö och lutar sig ut ur stigen.
En kille med vit skjorta spelar en vit gitarr.
En ung flicka visar sina vänner hur man använder en engångskamera.
En liten pojke som hoppar från en brygga ner i en sjö.
Damen med en grön mask på tandläkaren och hon ser väldigt olycklig ut.
En man med orange jacka och blå hatt som klättrar på ett snöigt berg.
En liten flicka med blont hår leker och plaskar i en lerpöl.
Ett barn cyklar nerför en gränd med graffiti i sig.
En gymnast bedöms vid ett tillfälle.
Folk går nerför gatan med en gatuförsäljare.
Mannen klädd i en traditionell klänning som klädsel, medan han står bredvid sin mula som också verkar vara klädd.
Två barn leker på en cykel.
Två män i motståndarlag spelar fotboll på ett fält.
En man hoppar och poserar för fotografer som ligger på marken.
Flickan tar en drink från en vattenfontän.
Spelunkern hittar vatten under sin vandring.
En man i en labbrock tittar genom ett mikroskop.
En blond tjej sover på en brun soffa.
En man sopar en trottoar utanför en tegelbyggnad under dagen.
Tre män lagar mat i ett kök.
En man på en ställning framför ett hus ler och poserar för fotografen.
Två tjejer i shorts håller hand vid en pool.
Fyra asiatiska barn sitter på en bänk och vinkar och ler mot kameran.
Barn cyklar i vad som verkar vara en utarmad nation.
En ung pojke, som bär kockmössa och förkläde, skär korv i ett kök.
Det här är en clown på en grundskola.
Den leende kaptenen håller i hjulet på sitt träskepp.
En gul bulldozer arbetar för att flytta smuts.
En kvinna i röd skjorta rider på en vit häst som galopperar längs träden.
En kvinna som sitter på en mycket stor sten och ler mot kameran med träd i bakgrunden.
Tre män i färgstarka kostymer tar sig ut på gatorna med peruker och galna solglasögon.
En flicka leker i en liten pool.
Två barn, en pojke i gul skjorta och en flicka i blå och vita ränder, svängande.
En man kastar ett fiskenät i viken.
En man med grå skjorta, blå jeans och neongrön skyddsväst står på en järnvägsbana med en vit lastbil och en vit byggnad i bakgrunden.
Två byggnadsarbetare lägger plåt över balkar.
Det finns ett band på scen med bandmedlemmar som bär inslag av blått.
En rockare med skjortan av sjunger in i en mikrofon medan han spelar trummor.
Jag ser en man som ställer sina saker från kundvagnen, redo att checkas ut.
Mannen med käppen är på en promenad.
En kvinna som bär vit skjorta fungerar på en ellipsmaskin.
En tjej som bär mask rider på en mans axlar genom en fullsatt trottoar.
Två flickor, en äldre och i svart och en yngre och i vitt, utför samma balettdrag framför dekorationer gjorda av ballonger.
Flera kvinnor utför en dans framför en byggnad.
En flintskallig man som går längs en trottoar medan han pratar på sin mobil.
En kvinna leker med fingerdockor som ett litet barn i en kostym går förbi.
En grupp människor ser unga män spela trummor med hjälp av provisoriska hinkar som instrument.
En tjej med normala och improviserade säkerhetsutrustningsrollblad.
En liten vit bil är på tågspåren och kan ha blivit påkörd av tåget bakom den.
Två rockare sjunger och spelar på en mörk scen.
En tjej med basebollmössa, vit t-shirt och blå shorts står i en berggrundsbelagd, skogsfodrad bergsström.
Två män som spelar gitarr inför en stor publik.
Ett antal människor dansar med sina betydelsefulla andra framför detta enorma hus.
Kvinna och hund säljer sina varor på den gamla byggnaden trappor utanför.
En kvinna och två män, som är klädda professionellt, har en diskussion.
En grupp män i röda och svarta jackor väntar på motorcyklar.
En kille klädd i vit uniform med nummer 3 på som spelar fotboll.
En man säljer snacks på ett sportevenemang.
Två män från det gröna laget tar itu med de andra medlemmarna från det svarta laget för bollen i en omgång rugby.
Barnen tävlar om att få tag i fotbollen.
En person i blått är den enda person som för närvarande kastar sin boll i en bowlinghall.
Flera fotbollsspelare på ett fält i aktion.
Ung man sitter på en skateboard, håller en mobiltelefon, och poserar på rulltrappan.
En kvinna klädd i blått som kör ett maraton.
Detta band gör sig redo att uppträda inför en publik i kyrkan.
8 för Iowa State stela armar en Texas AM spelare försöker tackla honom.
Två manliga curling spelare är på is sveper stigen framför polerad sten, en liten publik klockor.
Män spelar fotboll på ett lerigt fält.
En basketspelare i vita knäböj medan en spelare i rött rör sig mot honom.
Folk går genom en valvbåge i en gammaldags stad.
Två racerbilar, en röd och en blå, kör sida vid sida längs en racerbana medan de övervakas av flera åskådare.
En fotbollsspelare i vit uniform håller i en fotboll.
En mycket ung pojke stirrar framåt när han biter på ett litet föremål.
En kvinna och ett barn går nerför en gata.
En hockeymatch spelas med massor av människor som tittar på den.
Tre kvinnor studsar på bollar i gräset.
En afroamerikansk pojke med blå shorts, en svart och röd skjorta, och vita gympaskor, spelar tennis.
En man och en kvinna i vita skjortor kramar varandra.
En man som pratar med en familjeenhet som har någon sorts undersökningsapparat när de ser på och ler för att vara artiga.
Mycket ung pojke i en grön skjorta som ligger ansikte ner på en vit säng.
En extrem cyklist stannar för att vila när solen går ner i bakgrunden.
En kvinna skymmer i ett snöigt område och bär varma kläder.
Fyra flickor och en dam som lär sig att göra lite hantverk.
En man med svarta och vita ränder försöker stoppa en häst.
Herrn skannar bilden som kvinnan i den blå skjortan ger honom.
En kvinna med rött hår är hals djupt i molnigt blått vatten.
Två unga pojkar poserar med en valp för en familjebild.
Fyra barn tränar karate medan två vuxna tittar.
En mans lounger på en röd soffa i ett utställningsrum för möbler.
En grupp människor som pratar vid borden.
Två hästkapplöpning jockeys, en i rutig blå och röd och den andra i orange och brun, är racing mot en suddig bakgrund.
Den röda bilen ligger framför de två bilarna i bakgrunden.
En stor tjur siktar in sig på en man i en rodeo med sina horn, medan en rodeo clown springer för att hjälpa till.
En skjortlös man går mot en gul kajak.
En pojke på skjutbanan siktar och skjuter.
Två lag av pojkar som spelar fotboll i sanden.
Ett barn i blått och ett barn i vitt står på en kort betongvägg vid en bäck.
En kvinna ritar en blommig design på en lerkruka.
Folk går på en livlig gata i ett främmande land.
En högerhänt kanna för Saints kastar en pitch.
Två män, en i svart och vit och en i rött, spelar beachvolleyboll.
En man står i en båt och håller i lite nät.
En surfare som ramlade av sin surfbräda i havet medan han försökte rida en våg.
En tekniker som förbereder ett prov i labbet.
Fotbollsspelare hoppar i luften för att slå bollen med sina huvuden.
Två pojkar spelar fotboll mot varandra.
En äldre person går över en gata med ett paraply i händerna.
En grupp löpare springer mot två identiska skyskrapor.
En skateboardåkare rider upp en betongvägg och faller nästan av när han försöker ett trick.
Folk spelar ett spel i poolen.
En kille ger en kyss till en kille också
En man skriver en autograf i en ung pojkes bok.
En ung man i en blå skjorta slipar en räls på en skateboard i ett urbant område.
En asiatisk man sitter på spåret med lådor av jordnötter.
En brittisk gentleman, klädd i militäruniform, viftar med hatten med en bakgrund av människor som sitter tillbaka och tittar ut på vattenvägen.
Två bilar kör på en kapplöpningsbana.
En man i svartvit jersey håller gula skidstavar och förbereder sig för att lyfta.
Två människor lägger sig ner och kysser varandra på en gräsbevuxen gräsmatta.
Ett mycket litet barn i en denim baseball keps äter ett grönt äpple.
Fotbollsspelare springer för att få bollen.
En man i svart jacka och rutig hatt klädd i svarta och vita randiga byxor spelar en elektrisk gitarr på en scen med en sångare och en annan gitarrist i bakgrunden.
En man hoppar över en barriär från en tjur.
En kvinna i blå skjorta och vita shorts som spelar tennis.
En man spelar ett inlägg i en konsert
En man bär en stor massa metallbjälkar på axeln genom en skogsgård.
Kvinna med kamera kastar en frisbee för sin bruna hund att fånga.
Det finns en kontur av en man och en kvinna som observerar en brasa eller något annat stort brinnande träföremål.
Två flickor doppar händerna i en fontän när folk går förbi.
Ett vått, leende barn utan skjorta poserar med upplyfta armar.
Två män, den ene klädd i vitt och den andre blå, brottas.
En kvinna i en röd bikini som hoppar för att slå en boll medan hon spelar volleyboll på en strand.
Orange randig kattunge bitande blond flicka på näsan
En kvinna, som bär ett gult förkläde, tar av locket på en stor gryta.
Två barn korsar en liten bäck med hjälp av en stenbro.
Två afrikanerska kvinnor rider på en moped nerför en stad gata som verkar vara i ett väl överbelastat område i ett stort stadsområde.
Två pojkar framför en läskmaskin.
Cykelcyklisten bär svart, rider ner för en grusstig i en mountainbike.
En dam med tatueringar tar en bild av en målning med sin smartphone.
En kvinna i en mestadels svart outfit och vit hjälm rider en cykel med suddiga träd i bakgrunden.
Ett team cyklister rundar en krök medan närliggande åskådare hejar och fotograferar.
Fyra fotbollsspelare i svart är att ta itu med motståndarlagets spelare, visas i vitt, medan det regnar.
En löpare rusar efter yardage medan de förs ner av två angripare.
Basketspelaren i den vita uniformen med nummer 55 på vaktar spelaren i den svarta uniformen med nummer 10 på den.
En man pratar på en mobiltelefon utanför.
Professionella baseballspelare under All Star-spelet titta på en motståndare på fladdermus.
Smutsbiker gör en sluttande sväng i en skog under hösten.
3 basketspelare tävlar om bollen och en i röd tröja försöker ta bollen från killen i vit tröja.
En pojke tar tag i benet när han hoppar upp i luften.
Två barn som bär randiga tröjor och svarta byxor betslar utomhus nära ett spelset.
En man som bär solglasögon åker skoter.
En liten pojke som bär baseballregalia håller ett slagträ bakom huvudet med en baseball monterad framför sig.
Sex män sitter på ett fält av grödor som innehåller trälådor.
En brun hund plockar upp en kvist från en stenyta.
Det här är en man klädd i gult som håller i en brun hästs välde.
En man i vit skjorta och förkläde skär upp en fågel.
En latinamerikansk kvinna använder en wok utomhus för att laga mat.
Marathonlöpare tävlar på en stadsgata, med andra människor som står runt omkring.
Asiatisk kvinna bär solhat medan du cyklar.
En del barn är ute och leker i smutsen där det finns två träd.
En äldre man spelar ett arkadspel.
En flicka vid stranden av en strand med ett berg i fjärran.