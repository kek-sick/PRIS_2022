En grupp män lastar bomull på en lastbil
En man som sover i ett grönt rum på en soffa.
En pojke med hörlurar sitter på en kvinnas axlar.
Två män sätter upp en blå is fiskestuga på en is över sjön
En flintskallig man som bär en röd flytväst sitter i en liten båt.
En dam i en röd rock, som håller en blåaktig handväska som troligen är av asiatisk härkomst, hoppar från marken för en ögonblicksbild.
En brun hund springer efter den svarta hunden.
En ung pojke som bär en Giants jersey svänger ett basebollträ på en inkommande pitch.
En man i ett rörigt kontor använder telefonen
En leende kvinna i en persiko tank topp står håller en mountainbike
Ett litet barn står ensam på några taggiga klippor.
En person på en skoter i mitten av hoppet.
Tre små barn står runt en blå och vit tunna.
En kvinna sitter vid sin torkade blomsterutställning på en utomhusmarknad.
En kvinna som spelar en låt på sin fiol.
Tre personer på två smutscyklar och en fyrhjuling rider genom brunt gräs.
En halv naken man sover på sin stol utomhus.
En grupp människor som står framför en hydda på en parkeringsplats.
En ung kvinna gör mattor i regnskogen
Tre flickor gör ansikten när man tar en drink medan de står på en livlig gata.
En ensam man i svart t-shirt står ovanför publiken på en upptagen bar.
Kvinna och man går över trä rep bron med en varningsskylt bredvid den.
En man i kjol hoppar medan han jonglerar med knivar.
En asiatisk flicka i grön hatt och förkläde serverar drinkar på en bricka.
Byggarbetare som står ovanpå en maskin.
Två hundar leker med en orange leksak i högt gräs.
En söt bebis ler mot ett annat barn.
Tre män går på en väg i bergen.
En person parasailerar över en stor vattenförekomst.
En traktor rör på sig smuts för att hjälpa till att bygga upp en fasthållningsvägg.
En ung flicka som springer ensam i en park.
En person korsar gatan och undviker spill av färg.
Barn som leker på en lekplats, hängande på barer.
En person som bär en röd långärmad skjorta ligger på en vägg framför en lyktstolpe på ett mycket ovanligt sätt.
En grupp människor samlas runt en man i kostym och en liten pojke.
En kvinna sitter på en mörk bar.
Folk går nerför en trottoar där det finns en utomhusmarknad.
En man med en blå ryggsäck läser tidningen medan han väntar på att gå ombord på tunnelbanan.
En stor brun hund sticker ansiktet i sprinklern.
En blond pojke i en blå t-shirt står och ler inför ett hantverk av grönt nylontyg.
En ung vit hane sveper en veranda med en stor kvast.
En person som är mitt uppe i att kasta en grön bowlingboll nerför en bowlingbana.
Ett band spelar en rockshow för en barpublik.
En äldre man går en brun hund med rött koppel.
En man kör en gammaldags röd racerbil.
Unga vuxna bär röda, gula och svarta skjortor i en rak linje utför en skiss.
En ung pojke som kastar en sten i lugnt vatten.
Två kvinnor med kort hår är vända mot varandra och den blonda pratar.
En utstuderad figur står framför en ljust dekorerad byggnad.
En hund som går genom en liten bäck med en trasa i munnen.
Tre små hundar sniffar på något.
Två man paddlar kajak längs en flod med gröna träd på vardera sidan.
Två flickor går nerför gatan.
En grupp barn sitter i en skåpbil och tittar på en bok.
Beach goers tittar på ett hjärta kvar i himlen av en himmel författare.
När en flicka sitter lättvindigt på en offentlig plats, läser hon att hon håller boken öppen med handen som är en fjärilsring.
En man på en restaurang som äter lunch.
En man i kostym och glas har ett föremål i sina händer.
En man i svart våtdräkt surfar på en våg.
En kvinna med rosa handväska sitter på en bänk.
Tre kvinnor ler och sitter ner.
Ett rött plan som flyger över en båt när det spårar rosa rök.
En man i en sele klättrar på en stenvägg
Två byggnadsarbetare hjälper till med lastningen av en soptipp på en byggarbetsplats i städerna.
En kvinna i en färgstark outfit går förbi en vit lastbil fylld med flaskor.
En kvinna i blå hatt och gul kjol hoppar i ett område med syren.
En man bär gulddräkt medan han står med sin guldcykel.
Baby tittar på löven på en gren av ett träd.
En vaktmästare ska moppa på en tågstation.
Två små svarta pojkar leker med plastflaskor och har mycket kul.
Gröna trafiksignaler lyser upp när folk tittar på motorcyklar.
Två personer klättrar på en stenvägg med ett rep.
En man och en kvinna som fiskar på stranden.
Ett barn gör en backflip medan du hoppar på en studsmatta.
Barn rider en svängande karnevaltur
Två personer håller en stor upp och nedvänd jordglob, ca 4' i diameter, och ett barn verkar hoppa över Antarktis.
Två män i militären spelar baseball.
En kvinna i svart klänning kör en kärra med termos nerför en asfalterad gångväg.
En polis som stoppar ett fordon vid vägkanten.
Mannen står på en brygga bredvid en båt på en stilla sjö.
En grupp skotska officerare gör en demonstration.
En kvinna och ett barn sitter tillsammans i en dörrkarm längs en grå trottoar, när en man och två kvinnor går förbi.
En ensam brandman hjälper till att tämja en stor brand.
En person med lila skjorta målar en bild av en kvinna på en vit vägg.
En liten flicka ligger på golvet medan hennes yngre syster låtsas vara sjuksköterska.
En ung kvinna och äldre kvinna bär traditionell saris när de spinner textilier, tre personer är avbildade på bara midjan, och bär moderna kläder.
Kvinnor går genom djup snö och nerför en brant kulle.
FedEx-föraren lyssnar på arbetaren i den gröna hatten medan utrustningen lastas.
Den bruna hunden bär en svart krage.
En brun en vit hund springer nerför en gul och blå ramp.
Ett barn gör sig redo att läsa en bok.
En äldre japansk man som försöker fixa en liten röd och grå maskin.
Ett litet barn och en kvinna står runt en burd tupp.
Ett barn som är klädd som Spindelmannen ringer på.
En man klädd i brunt som håller i en lätt sabel.
En ung kvinna står och sjunger i en mikrofon medan en man bakom henne håller i en gitarr.
Två barn gräver hål i jorden.
Många av stolarna är tomma med bara ett fåtal människor njuter av solen.
En del män sitter på en båt nära en strand täckt av staplade stockar och pinnar.
En ung man bär något i en stor svart plastpåse.
En äldre, överviktig man kastar en pannkaka medan han gör frukost.
Män med gula kostymer står på scen med piano och en man spelar en upprätt bas.
Flera människor står nära träd vid skymningen.
En brun hund som tuggar på en stor träbit.
En vandrare poserar för ett foto i ett torrt fjälllandskap.
En grupp barn leker i vattnet under en bro.
En kvinna ler bredvid mannen som också ler medan hon håller i sockervaddkonen.
Två kvinnor står framför en klass av barn och pratar om en bok.
Två brunettkvinnor som pratar med ett klassrum fullt av blonda barn.
En person som bär hatt och halsduk ser åt höger.
Två personer går över en gata.
En gammal man håller upp en hund medan hans andra hund klättrar i hans knä.
Tre barn ser en man på scenen spela gitarr.
En pojke som tar en pinne från en flicka mitt i ett lopp.
En blå jeep kör ner i djupt, lerigt vatten.
Damen med svart hatt tar en bild medan snön faller.
En man som sitter på marken och spelar gitarr.
En hund trampar genom ett grunt vattenområde som ligger på en klippig bergssluttning.
En ung asiatisk kvinna hoppar mitt i luften i en trång stad.
Ett tremannaband uppträder på scenen.
Fyra personer protesterar mot Equinox behandling av unga arbetstagare.
En man som lagar hamburgare på en svart grill.
En man i en röd keps lutar sig mot en lätt stolpe.
En ung pojke i gul t-shirt hängande från en ring med andra barn runt.
Ett litet barn som äter frukt och dricker ett glas juice.
En man och två kvinnor i shorts, gå nerför gatan.
Två pudlar springer genom snön.
En rödhårig flicka bär en Spider-Man-dräkt medan hon rider en lekhäst.
Man i en liten vit båt på en sjö.
Skidåkarna är framför lodgen.
Folk fotograferas när de klättrar eller vandrar i bergen.
Flera personer simmar i en vattenförekomst.
Kvinnor i strand bikinin spelar volleyboll i det soliga vädret.
En man och en kvinna sitter mitt emot varandra vid ett restaurangbord.
En mor och två barn poserar med roliga ansikten.
En Golden Labrador simmar genom vattnet med en röd leksak i munnen.
Fyra män står nära en gul bil.
En grupp män, kvinnor och barn, alla klädda i hattar, pratar på stranden.
Lilla pojken i Cami kryper på brunt golv
En liten flicka donerar till Frälsningsarmén nära en butiksfront med vita plastbehållare.
En gul hund bär en boll i munnen på stranden.
En man i röd skjorta står med två fitlar framför en gammal struktur.
Mannen ser ut som en kvinna som pratar på en bar.
Ett band som spelar i en utomhusteater, längs floden.
Två kvinnor ler vid ett evenemang.
En kvinna i rosa skjorta som visar en man med randig tröja hur man gör lite arbete med garn.
Ett barn som sitter på en stenformation.
En man som sitter på en stol med en öl i händerna och steker något att äta på en träpinne.
En polis i uniform klädd i ett öronstycke.
Det finns en man i brandmannens utrustning som korsar vägen nära en vit buss och en röd halv.
En svart och vit hund som simmar i klart vatten.
Ett band spelar musik på scen på en konsert.
Det finns 3 personer som spelar musikinstrument och en annan person ser ut som hon sjunger.
En man som spelar tangentbord och sjunger in i en mikrofon.
En ung pojke hoppar ner i vattnet.
En kvinna läser ett kort medan hon sitter på en soffa, medan en annan kvinna står bredvid henne och håller ett glas att dricka.
Det finns byggnadsarbetare som arbetar hårt med ett projekt.
En man rakar sig medan han sitter på stranden framför havet.
En blondhårig kvinna som bär en blå skjorta packar upp en hatt.
Två män pratar med varandra bakom ett organ medan en ensam kvinna står till höger om dem.
En ung blondhårig man talar in i en mikrofon.
En betjänt på motell som bär en trenchcoat med en massa bagage.
Hund i växter hukar för att titta på kameran.
En grupp spelar musik på scenen inför en folkmassa.
Tre hundar leker i snön.
En man och en kvinna pratar medan de står bredvid ett träd.
En hund hoppar för en gul och svart boll.
En äldre dam i grå och röd tröja lagar mat.
Kvinnan i kappa utanför ett hus medan snön snöar
En kvinna som bär en annan kvinna i matchande träningskläder på ryggen.
Ett barn som står vid en barnvagn och håller ett leksakssvärd.
En kille med lockigt hår åker skateboard längs en grå ramp med gula bokstäver.
En man rullar ett cirkulärt bord tvärs över golvet.
En grupp människor sitter i en båt på en stor vattenförekomst.
En man i gul skjorta står på trottoaren och mäter.
En kvinna i blå skjorta och jeans kastar något i en container.
En kvinna i en dominomask och hårt hår är på fest.
En person parasails på krönet av en våg.
Män med blå uniformer sitter på en buss.
En ATV försöker ta sig ur ett dike.
En man tar itu med en annan man medan han spelar fotboll.
En fotbollsspelare i rött och vitt pratar med en tränare.
Två flickor sitter nära en vägg och tittar på ett sportevenemang.
En man som tränar för OU har solglasögon på huvudet under en fotbollsmatch.
Detta fotbollslag bär röda skjortor och röda hjälmar.
En pojke i svarta kläder gör ett hjul på stranden.
De poserar för en bild.
En man i grön skjorta kysser ett gråtande barn medan han tittar på löpare i en road race.
Fem medlemmar i ett band spelar en låt.
Tre kvinnor sitter på en filt på marken med ett barn, och pratar och har roligt.
En man och en pojke sitter vid ett altare båda håller klockor.
En man med solglasögon hjälper ett barn med solglasögon att glida ner för ett rutschkana.
En hund springer genom gräset mot kameran.
Flickan med lång hästsvans beredd att kasta bollen till en annan spelare på fältet.
Två män brottas på gult och blått golv.
En tjej i röd och vit skjorta och blå shorts gör sig redo att kasta en boll.
En sittande man arbetar med sina händer.
En brun hund springer på sanden med en käpp.
En person roddar i sin båt i vattnet.
En man i röda och vita randiga skjortor sitter på en pall vid ett korvstånd.
En man fotograferar vita och gula tulpaner.
Två män på Fez har en diskussion på en utomhusmarknad.
Man och pojke leker med hund vid solnedgången på en strand.
En varmluftsballong som rör sig ner med en mans skugga i bakgrunden.
Den här mannen bär en vit keps eller hatt.
En kvinna som får en ansiktstatuering av svarta linjer och glitter.
Ett litet barn i en denim hattar spelar i ett däck.
En skara människor står på gatan framför en serie vita tält.
En massa människor går genom parken.
En mörkhårig kvinna med blå blus och solglasögon håller en banderoll medan en ung flicka med flätat hår skriver på banderollen.
Många asiatiska barn gjorde ett tåg under ett viet namtecken.
En cowboy vred en häst i en rodeo som hästen gör en ryggspark
En brud och en brudgum på deras bröllop kysser
Två räddningsarbetare lägger block under ett tåg.
En man som jobbar på järnvägen på en järnvägsstation.
Vissa byggnadsarbetare, det finns betong som blandas i skottkärror, de bygger eller reparerar en vägg, väggen är fortfarande våt.
Ett band som spelar på trottoaren.
Män i orange kostymer tittar på en maskin gräva nära vad som ser ut att vara tunnelbanespår.
Unga vuxna som klär sig lättvindigt går omkring på ett fält.
Den stora bruna hunden rinner genom grunt vatten.
En man och kvinna går över en tom gata.
En man i det kalla vädret i en hink som arbetar på en kraftledning.
Två barn i gula jackor leker i lera.
Det finns flera personer som går över en slinga på en inverterad berg-och dalbana.
En kvinna och en liten pojke delar en stol.
En grupp människor står i en lös linje på en tegelmark.
En ung flicka simmar i en pool.
En pojke med orange skjorta ler, medan en pojke i blå skjorta ser på.
En liten flicka står i en pöl utanför.
En liten blond tjej håller i en smörgås.
4 personer försöker fixa en cykel på en park
En mycket våt brun hund växer fram ur vattnet.
En hund springer över ett fält med en boll i munnen.
En grupp människor väntar bakom en barrikad och ser åt höger.
Ett barn som bär en röd tröja hänger upp och ner från ett träd.
En karnevalspelsoperatör tar pengarna från två villiga tävlande.
En pojke ler för kameran i en grupp sittande barn.
Två barn utan skjortor sitter på kanten av en fontän.
En man drar på sig tröjan när en kajak lägger sig vid fötterna.
En gammal man som går med en mapp i handen
En ointresserad ung kvinna och en äldre man står vid en bar.
En ung blond pojke hoppar från sängen till sängen.
Ett litet barn svänger tillbaka ett rött basebollträ.
Han pratar på mobilen framför en sportaffär.
Här är två mammor som lyssnar på ett litet barn.
En kvinna i blå skjorta spelar ett instrument.
Detta är en fullsatt korsning i en stor stad på natten.
En man som sitter i klart grunt vatten vid en stor klippa.
Ett par vandrare tar en paus för att ta en bild.
Fyra goth ser människor som går nerför en gata med träd i bakgrunden
4 personer är fastspända vid en nöjespark rida
En pojke gör ett skateboard trick från en metallplanka.
En man på en strand som bygger ett sandslott.
Den stora bruna hunden jagar den lilla bruna hunden.
Män i vita kläder håller upp sina händer.
En kvinna thows en frisbee till en hund som en baseballspelare i uniform kör bakom henne.
En svart hund som står i något gräs och håller ett vitt plastföremål i munnen.
En båt med människor och deras tillhörigheter ligger i vattnet.
Ett paket cykel road racers lutar genom en kurva.
Tre personer sitter utanför vid ett bord med konstverk som lutar sig mot det.
En vit kvinna och svart man som går nerför gatan.
En man i en vit t-shirt målning mitt på en stenlagd väg.
En brun, svart och vit hund som skäller upp ett träd.
En man i blått och rött ansikte målar för en bild med en kvinna.
Två pojkar spelar ett spel med kulor.
Två män väntar i baksätet på en bil medan föraren går in i förarsätet.
En pojke rider en sväng.
En svart man tittar på en annan svart man som leker i vattenfallet.
Person med en röd backpackers går på en vandring.
En asiatisk frukt- och grönsaksförsäljares urval av bananer, apelsiner, meloner och mycket mer i sin lilla båt.
En stor publik står och tittar på med en stor byggnad i bakgrunden.
Tre kvinnor i mörka sjalar och hattar pratar på en tegelgata medan en hund sitter bredvid dem.
En man i vit skjorta gör shish kabob.
En person med neonrosa hår och gul skjorta tittar ut över en strand.
Man tittar på en kvinna som röker på trottoaren.
En man i svart skjorta och bruna lastbyxor som håller en spade ovanför huvudet.
En man som slickar ansiktet på en kvinna i glasögon.
Det ena barnet går före det andra.
Den unga flickan får kaninöron av den unge pojken bakom sig.
En ung baby, klädd i rosa fleece outfit, ler medan den ligger på höstlöv.
En närbild av en kvinna med kort rött hår.
En fotbollslagsspelare i en grön skjorta springer iväg från fältet.
En flicka leder sin hund över ett hinder.
Flera barn höjer händerna medan de sitter på en färgglad matta i ett klassrum.
Sailors står på toppen av en gangplank till en stor båt.
En medelstor vit hund hoppar upp för att fånga en liten duk Frisbee.
En man i grå t-shirt vilar.
En svart hund hoppar genom vatten och håller en käpp i munnen.
Två svarta hundar som springer ner på vardera sidan av en asfalterad väg
Fyra personer i tillfälliga kläder står utanför och håller soppåsar.
Folk och kameler tar en paus i öknen.
Fyra hundar leker i en cirkel och en svart hund går sin väg.
En man i en arméuniform talar in i en mikrofon.
En grupp asiatiska människor på en autoshow stirrar och tar bilder på ett nytt fordon.
En simmare som simmar i en simbassäng.
Kvinnan med en vit skjorta och bankerna ligger på en soffa inne i ett hus.
En man sänder handsignaler bredvid två unga flickor.
Tjej i vit skjorta blåser bubblor i mörkt rum.
Pojkar och flickor från en östlig nation som ler på ett fält.
Ett barn i orange skjorta hoppar av balar av hö medan andra barn tittar.
Pojke gör tricks på en skateboard
En man sträcker sig upp för att arbeta med kablar ovanför ett skrivbord.
Ett litet barn sitter vid ett bord och äter ett mellanmål.
Fyra barn som bär ryggsäckar vänder sig mot kameran och ler när de går på en landsväg.
En man med dreadlocks kopplar sitt öra för att höra ett telefonsamtal.
Mjuka stora skivor staplas på en spindel i en industriell miljö av en man när en annan ser på.
En hund på ett gräsfält som tittar upp.
En kvinna och ett litet barn har kul när de spelar brädspel.
4 barn sitter på en avsats och samtalar.
Den lilla bruna hunden är mitt i krukväxterna och fällda blad.
Två män målar en byggnad medan en tredjedel går förbi på sin mobil.
Vissa män tittar på en datorskärm på ett kontor.
Två kvinnor undersöker ett foto på en kamera.
En blond kvinna i en brun cowboyhatt gör en obscen gest mot kameran.
Den vita och bruna hunden springer över gräset.
En tonåring som läser en bok i klassen med anteckningar på skrivbordet ser uttråkad ut.
Två små flickor går längs löven.
En brud justerar sina män blomma på hans rock när hon håller sin egen bukett av blommor.
Kvinnan placerar en apelsinros som en boutonniere på mannens klädkrage.
Två kvinnor med sina barnvagnar som går längs en lövtäckt gata.
Fyra kvinnor klädda i roliga kostymer.
Denna gamla asiatiska kvinna vilar och beundrar sig själv på en till synes het dag i staden.
Tjejer i svarta bikinis som spelar beachvolleyboll.
En man med glasögon och en liten flicka med flytväst som simmar i en pool.
Tre barn bär bruna skjortor och jeans hoppar utomhus med löv på marken.
En kvinna fokuserar på sitt curlingspel.
En person bär många väskor.
Ett barn nära en blå scen med en färgstark varelse på sig.
En pojke står fånigt mitt i en social sammankomst.
Detta barn är i ett klassrum, klar för dagen, kanske
En man Wakeboards i vattnet.
Barn stirrar ut genom fönstret i en blå byggnad med röda fönsterluckor.
En salt-och-pepper-hårig man med skägg och glasögon bär svart sitter på gräset.
En kvinna och hennes två barn är på stranden och kvinnan hoppar högt upp i luften.
Ett par män som går på en allmän stadsgata.
En kille gör ett cykeltrick i en park.
En man i en färgstark skidjacka står med andra på en europeisk gata.
En kvinna i gul t-shirt och solglasögon går nerför en trottoar.
Två kvinnor ser ut över många hus nedanför.
Två stora hundar frolic i ett gräsfält.
Folket är klädda i tunga kläder och rör sig tillsammans.
En grupp människor som äter på en restaurang.
En kvinna som bär en svart t-shirt verkar gå upp i en rulltrappa.
Ett rum fullt av sittande och stående vuxna och barn, och åtta rosa och svarta ballonger hängande från taket.
En man och en kvinna poserar tillsammans på en kullerstensgata.
Två hundar springer och leker i snön
En liten hund som hoppar på en gata.
En man som bär en svart t-shirt spelar sju string bas en scen.
En pojke och en gammal man med käpp pratar.
En tjej med vit skjorta, svarta shorts och ett pannband spelar volleyboll.
Två män står på gatan täckta av graffiti.
En pojke i t-shirt och shorts håller i en snöboll och vänder sig mot ett snöigt berg.
En människa hänger glidande i havet.
Två husarer sitter upphängda på hästar, klädda i extravaganta ceremoniella kläder, var och en håller en sabre i sin högra hand, regerar till hästen på sin vänstra.
En hund som springer genom djupt snötäcke.
En medelstor grupp människor poserar framför kameran.
Stor brun och vit prickig hund som ligger på en jacka på gatan.
Två tonårsflickor har ett kort som hänvisar till perioder när de ler.
En mor och en son som ler när de slädar utför.
En man i svart skjorta kokar ur en kokbok i ett rörigt kök.
En kvinna i vitt spelar en svart gitarr.
En snowboardåkare hoppar i luften bredvid skidliften.
Flera personer står i ett rum och äter.
En man i hatt spelar ett ovanligt instrument för kontanter bredvid tunnelbaneutgången.
En kille maler en fönsterbräda nära en gammal väderkvarn
En kvinna i vit skjorta och svarta byxor hula hoops som en stor grupp människor ser på.
En äldre man intervjuar en annan i en tävlingsdräkt.
Två män i röda dräkter som utför kampsporter.
Ett litet barn rider en motorcykel genom leran.
Ett barn som bär hatt och jacka springer utomhus på en stenyta.
Ett barn som sitter på sin pappas axlar i en folkmassa.
Två gamla män i hattar slumrar i solen utanför.
Två pojkar i ett tält ler mot kameran.
En varmklädd kvinna i svart knäböjer med en liten brun hund nära en skara åskådare.
Två män sätter upp en elektronisk utrustning.
En kvinna som bär på en handlare Joes väska har somnat på tåget.
En bicyklist gör ett trick i luften.
En ung man i en grön tröja läser en tidning på stranden.
En man i grön jacka ler.
En man klättrar uppför en brant bergvägg med en säkerhetssele på
En ung man rider en självbyggd cykel tvärs över gatan.
Två bruna hundar brottas på den gräsbevuxna kullen.
Person i en lång röd rock som går framför en byggnad.
En utländsk kvinna sitter med mycket färgstarkt tyg.
Två pojkar i ett stängsel hoppar i luften medan de håller i en basketboll.
En man med glasögon i mikrofonen tittar ner på papper i handen.
Ett barn med grön skjorta håller en röd boll mot munnen.
En man med en tatuering på armen som lagar något i en stekpanna.
Ett band på fyra som spelar ett gig.
En grupp unga asiatiska män som går i maraton.
En man som drar föremål på en vagn.
Tre stora hundar njuter av en romp i snön.
En fågel flyger över vattnet.
En grupp föräldrar sitter vid en utomhussammankomst.
En gul bil går snabbt längs ett snöigt fält.
En grupp barn satt och spelade sina instrument.
Grupp av vuxna som sitter runt bordet och lyssnar på presentationen
En kvinna klädd i grön skjorta läser av en projektor för sin klass.
Ungdomar är engagerade i ett spel.
Bollspelare i blå och vita uniformer är på planen och spelar baseball.
En kvinna och två pojkar tittar på en informationsstation.
En grupp människor som driver ett välgörenhetsmaraton.
Två kvinnor står med skidstavar i djup snö.
Alla står tillsammans framför en staty av ett djur, och de bär alla coola kläder.
En ung skidåkare tittar på kameran.
Två unga flickor klädda i rosa pyjamas sitter på golvet framför stora fönster som leker hus.
En kvinna och barn rider kameler nära havet.
En man ler med en hand i pannan på en fullsatt bar.
Gatan är full av folk med kappor på.
Två män i ett främmande land ler, en står och en sitter med korsade ben.
En liten brun hund springer på gräset.
En nattlig gatuscen av en restaurang.
En snowboardåkare gör ett trick.
Asiatisk kvinna i postförsändelse uniform driver en stor hög med paket.
En kvinna i blå skjorta cyklar.
En kvinna i vit tennis outfit hoppar upp för att träffa bollen.
En ung kvinna övar ett stränginstrument inomhus.
En brud och brudgum tar bilder medan två män står i närheten.
En kvinna som håller en vit och svart hund.
En pojke i röd skjorta som försöker spela gitarr.
En ung expedit som letar efter nya mejl från kunder.
Tre äldre kvinnor i ett vardagsrum, dekorerade för jul, en "VAIO" anteckningsbok är centrum för uppmärksamhet.
En vit fluffig hund hoppar och fångar en leksak.
En matador i en färgstark outfit rider en tjur
Barn badar i vatten från stora trummor.
En brun och vit hund hoppar upp med en gul boll i munnen.
En grupp människor i blå skjortor på ett sportevenemang.
Tennisspelaren bär en gul och blå skjorta och ett blått pannband.
Två små flickor i blå klänningar skrattar.
En liten flicka i en rosa tutu övar dans med halsdukar.
Två personer springer på toppen av ett berg.
En grupp kvinnor dansar Bali stil i färgglada kläder och makeup.
En cyklist som hoppar i skogen.
Flera människor går bredvid ett vitt staket i ett främmande land.
Kvinnan står på en tegelvägg och tar en bild
En kvinna som bär vita shorts, gula topp och vita sandaler verkar kasta en pinne.
En person kör sin smutscykel.
En liten flicka av asiatisk härkomst, sitter i en svart hink och äter en marshmallow, med ett stort leende i ansiktet.
Två terrier leker på trägolvet i sitt hem.
En liten pojke med napp och en röd skjorta leker med en trädgårdsslang.
En tonårspojke på en cykel gör tricks.
En gammal man i svart jacka tittar på bordet
Mannen i den blå skjortan går med mannen i rött.
En kvinna som hänger i ett träd, hennes ben inlindat i tyg.
En ung barfotaflicka som bär hjälm går nerför ett mossigt täckt fallet träd.
En svart hund hoppar över en mångfärgad barriär.
En pojke i blått, spelar fotboll, på väg att sparka bollen.
En besättning av cykelmedlem gör sig redo för ett lopp.
En kille flyr från en svart tjur.
En pojke med en mohawk som jagar gäss i en park.
Liten brun och vit hund som springer på trottoaren.
Två barn sätter sina ansikten i en riddare och kunglig kvinnas bild.
Skuggan av två män på riggning.
En svart pudel leker med en annan hund i ett torrt fält.
Flera människor njuter av en cigarett nära ett askfat.
En vit hund med bruna märken hoppar ner från stranden i vattnet.
En fotograf tar ett foto av ett meddelande på en uppsättning dörrar.
En liten flicka i en rutig klänning leker med sin stora blå boll nära ett mesh staket.
En man tränar boxning
En grupp ungdomar poserar i luften på en sandstrand.
Kvinnan håller i en fiol.
Resenärer på en mycket kall dag vandring.
En man i grå skjorta gör ett skateboardtrick i trappor.
Tre män går bredvid ett tält med en skylt på.
En ung flicka som står på ett gräsfält.
En pojke i grön och gul klänning lär sig boxning.
En man och en kvinna som leker utanför.
En ung flicka som bär klänning och sandaler springer i gräset.
En kvinna med lila hår och en man i militära regalier.
Folk dansar och klappar där med händerna.
En man stirrar på ett förbipasserande par när han går nerför kvarteret.
Mannen i vit skjorta och randiga shorts spelar organ observeras av människan bär gul skjorta
En stor grupp människor tittar på en artist på en scen.
Bilen lämnar ett dammspår när den går runt grusspåret.
En grupp människor lyssnar på en man som pratar utanför.
En skäggig skallig man i en solbränd randig skjorta vilar huvudet på en annan mans arm.
En pojke förbereder sig för att sparka ett mål skott
En cykelcyklist cyklar på vägen bredvid klippor med snö.
En långhårig post svänger runt hans våta hår i havet.
En pojke och en man klädd som rodeo clowner stående i sand
En ung flicka ler och sticker tummen upp medan hon poserar framför en sköldpadda.
En man i blått cyklar på ett spår.
En enda person fallskärmar genom en lugn solnedgång.
En servitris står bakom en disk full av kakor.
Två cyklister korsar gatan på en mycket breezy Kalifornien dag.
En grupp musiker spelar in musik.
Två personer spelar vattenvolleyboll i en pool.
Det finns ett café i ett gathörn med en oval målning i hörnet av byggnaden.
En pojke lyfter upp en annan pojke på ryggen.
En kvinna som använder en stor kamera medan hon står på gatan.
En flicka bär en stor blå och röd hatt.
En kvinna applicerar ansiktsfärg medan en pojke med en Mohawk håller i en spegel.
Flerkulturell grupp vuxna på en samling, en man med tatueringar kastar något.
En man i blå skjorta rider en enhjuling med flammande batonger i handen.
Ett litet barn leker i en vattenspridare.
Fyra barn leker på verandan medan deras far tittar på.
En man håller ett spädbarn medan han lutar sig mot en byggnad.
En kvinna med två medaljer runt halsen som håller upp sju fingrar.
Männen slåss under matchen.
Två flickor äter tårta och en har blå glasyr i ansiktet.
En kvinna sätter en hjälm på en liten flicka.
En publik är utanför och tittar på någon i mitten av dem.
En pojke i en park som leker med två apelsinbollar.
En ung blond flicka som står på en kudde på en säng och ler med slutna ögon.
En man sjunger in i en mikrofon medan han håller i en gitarr.
Man med Mardi Gras Pärlor runt halsen håller stången med banderoller
En man i grönt och en kvinna i svart stretching.
En man tar ett foto av en annan man och hans två hundar på några gräsbevuxna kullar
En man som gör en offentlig show med eld.
En stor svart hund springer längs ett staket i gräset.
En motocross ryttare är något luftburen på en tävling kretshopp.
Det finns en kvinna som cyklar nerför vägen, och hon knäppte en wheelie.
Den svarta hunden hoppar över vattnet mot en frisbee som flyter nära en båt.
En man i svart jacka och svart hatt spelar trumpet.
En man klädd i grön snowboard på en bänk.
En indisk man sitter utanför en restaurang vid ett bord.
Tre män i kostym sätter ihop händerna.
Små hundar i kostym står på bakben för att nå dinglande blommor.
Man glider ner för trappan ledstänger på en cykel.
En man med en hink och en flicka i hatt på stranden.
Folk går på en trottoar framför en bar och grill.
En stor hund hoppar i en fontän medan en man i svart T-shirt och väst står i närheten.
En man på en båt med orange byxor som håller i ett rep.
Två män är ute på en ljus, solig dag och försöker fånga lite fisk på sjön.
En man står på byggnadsställningar och målar en vägg i korallfärg.
En försäljare sitter mitt i en uppvisning av glasögon på en gatumarknad i ett asiatiskt land.
Två personer med vita skjortor som går uppför trottoaren och pratar i telefon.
Den lilla flickan med det gröna halsbandet springer iväg från nätet.
En konstnär målar utanför.
Två asiatiska barn, en pojke och en flicka, står på golvet bredvid ett träd.
Folk i kö gör sig redo att gå ombord på en buss.
Två lag, ett i rosa och ett i vitt, spelar lacrosse på ett fält.
En kvinna som bär en gul hjälm använder en zipline.
En svart hund som simmar i vattnet med en tennisboll i munnen
Tre män rider i en mörkblå bil.
Med ett badkar som vilar på yttertaket, flaggor fastsatta, är bilen redo att lyfta för rallyt.
En man i blå skjorta som blåser i en trumpet.
En manlig metallarbetare som använder ett svetsverktyg i sin högra hand, medan han håller masken i sin vänstra hand, i ett mellanlägset eller lägre klass område.
Många står vid en fontän under ett blått och vitt paraply.
Kvinnan syr för att försörja sig i sitt land.
Gatuförsäljaren rätar ut varor på bordet.
Tre män står runt en vagn nära några motorcyklar.
En bankkassor står vid en disk.
En man i röd luva med ett vitt förkläde står framför en väggmålning.
En man tittar på en av sina fyra plattskärmsdatorer.
Två människor rider sina cyklar på en grusväg
En ung smutsig asiatisk flicka som bär på en kudde.
Ett barn som är på stranden av en sjö som pekar ut något i himlen.
Ett par äldre pojkar spelar gitarr.
En man i vit skjorta och khakibyxor hukar sig på en fallen trädstam.
Två pojkar förbereder en liten segelbåt när två flickor tittar på dem från stranden.
En gammal man klädd i sjukkläder håller i en yxa medan han står på en kulle.
Tre personer är på stranden och knäböjer eller står nära vattnet.
En man i en gul topp står framför ett litet skjul, sett ovanifrån genom trådnät.
Ett barn är motvilligt på väg att bita i en svamp.
Två kvinnor bär rosa T-shirts och blå jeans konversera utanför klädaffären.
En uppsatt polis på en fallfärdig häst undersöker en folkmassa.
En stor svart hund gräver i den djupa snön.
En man fotograferar en sjö med berg i bakgrunden.
En brunettkvinna i ett Robins äggblått förkläde mjölkar ett brunt djur.
Folk protesterar mot åldersdiskriminering i ett organiserat gatumöte.
Två unga flickor spelar basket, en i vitt försöker lägga sig medan den andra i rött försvarar.
En kvinna i bikini som gör ett hjul i sanden.
En man med brun skjorta, grå väst och svart keps spelar elbas.
En kvinna med blont hår dricker ur ett glas.
En ung pojke som låg på en sjukhussäng med benet över sidan.
Två medelålders män i ett rum med musikutrustning talar med varandra.
En hunds mun öppnar sig för att avslöja sina skarpa tänder.
En äldre indian man och kvinna i deras hem.
En man lägger sig på en snöbank som har staplats högt runt ytterdörren till sitt hus.
En ung flicka sträcker sig ut för att klappa en hjort.
En kvinna med svart hår, klädd i svart topp och röd kjol skakar näven mot någon.
En man som knuffas i rullstol genom ett bibliotek.
Två hundar ligger i snön med munnen öppen.
En vänligt inställd kvinna städar golvet i sitt vardagsrum.
Två hockeyspelare redo att starta spelet med domaren av dem på väg att släppa pucken.
Runners passerar en kontrollstation i staden.
Grupp av människor som dansar på en klubb eller fest i kostym.
Två barn förbereder sig för en elefanttur.
En ung vuxen som bär jeans och en kamouflagetröja som spelar en svart elgitarr.
En person klädd i en gul animerad dräkt i ett offentligt område.
Simmare i en sjö som bevakas av en pojke som sitter på en vägg.
En skara människor på en stadsfestival med rök och fyrverkerier
Hund på koppel hålor i snö på landsbygden.
En grupp läger i ett öde område.
En kassörska med en svart god tröja räknar växel.
En pojke som får håret avspikat av sig av en annan pojke.
Här är en bild på en tonåring som klipper sin brors huvudhår.
Turisten tog bilder på en byggnad i Kina.
Pottery och bilar visas på en parkeringsplats med en man i en blå outfit lutar mot framsidan av sin bil.
Två män bakom en cirkulär bar i ett rum fyllt med människor.
Män och kvinnor väntar på att tåget ska stanna.
Barnen samtalar och lär sig i klassen.
En man sjunger in i en mikrofon medan hans band spelar.
En sångare uppträder tillsammans med publiken.
En äldre kvinna som bär blå hatt sitter på trottoaren och hugger något gult på en bräda bredvid henne.
En byggnadsarbetare i svart skjorta och jeans sätter upp sin stege.
En servitris i en vit t-shirt som serverar gäster på en restaurang.
Blondhårig man klädd i en svart fleece jacka skulptering.
En tjej som tävlar i gymnastik utför en modig rutin när hon imponerar på publiken.
En konstnär som arbetar med en isskulptur
En man i blå rock drivs på sin släde av två hundar.
Det här är något slags band eller symfoni som övar.
Två personer spelar ett spel mot varandra.
Flera flickor leker med mjöl.
En ung flicka spelar ett musikinstrument och sjunger in i en mikrofon.
En man som spelar Mike Tysons Punchout på sin dator.
En man som ser ut att ha blivit träffad ligger på marken framför något skräp.
Scen av en person som skyfflar snö medborgare som går runt i en kall vinter miljö
En grupp människor i rutiga kjolar, svarta västar och vitkollade skjortor spelar trummor.
En kvinnlig konståkare i en röd jacka övar sina rörelser.
En grupp människor som springer ett maraton på vintern.
En kvinna och en pojke på scenen skrattar med ett tält i bakgrunden.
En svart man i kockrock är i telefon medan två andra män i förkläden skrattar.
En ung flicka som går längs sidan en liten bäck
En brunettkille i en brun blazer pratar med en publik på en komiker show.
Två barn som dansar på en dansuppvisning.
Här är en bild på en kvinna och hennes man och barn som tar en promenad vid parkeringen.
Lynyrd Skynyrd uppträder på en konsert.
En man och en kvinna sitter på en bänk och ser en båt gå förbi.
En stadsgata har många tecken på kinesiska.
Flera personer pratar och tillbringar tid tillsammans i ett rum.
En grupp musiker som spelar musik på gatan.
Den här mannen verkar försöka göra något slags politiskt uttalande i en upptagen stad.
Två barn som leker på ett djungelgym.
En man sitter på dörrtrappor framför ett hus.
En man i kostym går på en livlig gata.
En man i vitt förkläde och hatt säljer kött på en livlig gata.
En kvinna står och bär en grön och gul halsduk.
En äldre asiatisk kvinna bär en beret, solglasögon, en gul halsduk och en rutig jacka.
Människor sitter bland vissa pelare medan en annan person går förbi.
En man och kvinna veterinär kollar en mycket stor tiger som ligger på marken.
Två personer tittar på kläder i ett skyltfönster.
En man med ryggsäck sitter på en grusväg och pekar mot horisonten.
Två män sitter runt en skinande grill.
En kvinna i gul jacka som följer två andra kvinnor.
En man i rock pratar på sin telefon på gatan.
En pojke bär en grön skjorta på en cykel som reflekterar från ett skyltfönster.
En liten flicka som kikar över en blå vägg.
En ung man får något att äta i en munkkoncession.
En gammal man sitter med en bricka i knät.
En afroamerikansk man i solbränd hatt, kostym och solglasögon står vid en tegelvägg.
Tre män pratar framför gamla trappor på gatan.
Svarta är i mataffären för att komma dit med mat.
En man och två barn som korsar en gata.
En man i kostym som röker cigarr och läser en tidning som går på gatan.
En grupp människor som spelar gitarr i vitt.
En hund hoppar i luften för att fånga en apelsinfrisbee.
Flera personer står på en tunnelbaneplattform.
De tre barnen är i en bur.
Två personer står framför en byggnad.
En äldre kvinna som använder ett rosa paraply för att skugga sig från solen.
En baseballspelare sparkar upp smuts som glider framför en fångare.
Två kvinnor i blå kostymer sitter på cementen utomhus med betong och långa glasfönster bakom sig.
Två män som röker utanför en park.
En man i blå skjorta har ett tecken som säger: "Kom igen nu, vad är gayare än te."
En kvinna i grön skjorta går nerför en fullsatt gata.
Två kvinnor som sitter i silverstolar och väntar på tåg eller tunnelbana i en inomhusstation.
En folkmassorna i närheten av början av ett maraton.
En ung pojke bär en grön, vit och röd flagga och går bredvid en kvinna.
Många människor samlas för att titta på två män som är ett instrument och håller ett tecken.
En man i en svart och vit randig skjorta som fotograferar en kvinna vid en fontän.
Två personer sitter på en cementbänk och chattar över lunchen.
En militär man som håller i en kamera och visar ett barn filmen på kameran.
En man knuffar stolar på en livlig gata.
En man som håller i en mikrofon och pratar med en grupp människor utanför.
Två män samtalar nära en vägg med graffiti på den.
En tjej med ansiktsfärg och en orange tröja står med sin fest.
En person står bredvid ett trästaket med blommande träd i närheten.
En vältränad ung kvinna kickboxar med en röd boxningssäck på ett gym.
Lemonade ståthållare arbetare sätta upp butik för dagen.
En man sitter i ljust färgad grön och blå monter med annonser bakom sig på gatan.
En ungdomsfotbollsmatch där tre ungdomar kämpar för en fotboll.
En man håller ett barn på sina axlar när ett folk går runt honom.
En man i ett förkläde som står framför maten under en meny.
Street scen av blond kvinna i guld rock och rosa mini-kjol framför en bakåtvänd polis motorcykel.
Flera artister klädda i vita kläder och maroon hattar är uppradade mot varandra.
En vit blond dam som bär en blå väska och åker skoter.
En kvinna som sitter på en offentlig bänk.
En grupp människor sitter vid ett bord utanför och dricker och pratar.
En liten asiatisk flicka springer in i fokus på en tegelgata.
En kvinna och fyra barn korsar en livlig gata.
Kvinnor i etniska kläder sjunger tillsammans.
En kvinna pratar med en ung flicka över en disk.
En kvinna grillar god mat i parken.
Polisen brottas med en man med handen uppe i luften när andra poliser tittar på.
En man i svart skjorta sjunger in i en mikrofon.
Två unga män i blå jeans och sneakers korsar en stadsgata.
Två tjejer leker på ett träd med sin hund.
Det finns en ung kvinna med en väska som ler framför en byggnad.
En man och en kvinna går nerför en stig vid vattnet mot en hängbro.
Tre kvinnor springer barfota på sanden mot vattnet.
En bebis som sitter på en blå cabriolet.
Två män tittar på skärmen på en bärbar dator medan en typ och en poäng på skärmen.
En färgstark parad ledd av en man som bar en röd flagga.
En man i grå hatt och tank topp med svarta shorts gör en handstand.
Kvinnorna håller pojken medan de tittar tvärs över gatan.
Bilden visar återspeglingen av en man och kvinna som befinner sig vid en terminal av något slag.
En man plockar upp en drypande kvinna lyckligt.
Mannen i det vita bältet och solglasögonen håller flickans hand.
En man går längs trottoaren bredvid en gata.
En man som bär olivdrabbkläder håller sig upp från marken med händerna.
Fotografer på en plats som gör en dokumentär.
Man och kvinna i svart står nära varandra på gatan.
Folk som deltar i en J.P. Morgan Corporate Challenge.
Flickan och pojken kysser varandra medan de sitter på en träbänk.
En man som bär glasögon går ut genom en pool vid stegen.
Det finns en ung kvinna klädd i grönt och rött med en mexikansk flagga ansiktsmålad på kinden.
En hjälmcyklist som flyger från en ramp i skogen.
Två kvinnor klädda i vitt och med höga klackar går på gatan.
En indisk man går förbi ett tempel på sin väg för att be.
En välbyggd svart man står i tunnelbanan och lyssnar på hörlurar.
Två män sitter utanför och pratar med ett gratisrådstecken.
En kvinna i röd klänning med rött hår som står framför ett ljust, flerfärgat hem.
En kvinna är rullskridskor i en skum uniform.
En kvinna i svart klänning och fluffiga öronmuffar som går nerför gatan.
Det finns många människor i en byggnad med en del människor som lagar mat.
Folk provsmakar mat från ett bageri på en lokal potluck.
En utsikt över en gata kantad av stora, rena byggnader.
En flicka med blå dreadlocks sitter på vägkanten.
En man i Denver Broncos jersey är med sina vänner.
En kvinna som blir underhållen av en clown på en lokal mässa.
En man i en lång blå mantel går in i en gammal stenbyggnad.
En dam i en ljusrosa skjorta drar en varm matvagn.
En person med långt blått hår som står bakom en stor skara människor.
En grupp strandbesökare håller i händerna och bildar en linje mot vattnet, nerför stranden.
En man i vit skjorta spelar fiol på gatorna.
Många går på en grusväg och har sommarkläder på en solig dag.
Två personer i helkropp solid färg spandex kostymer sitter i stolar i en publik.
En svart man med mössa sitter i en buss.
En gentleman som kommer ut ur en tvättomat.
En man i kostym och slips i en tjusig byggnad pratar på podiet.
Mannen har somnat på soffan.
Fem män som alla bär vita rockar står bredvid lamm i ett slutet område
Två vattenskotrar, en röd och en vit, gör ett stort stänk i vattnet.
En grupp på fyra personer fotograferas från en bil.
Folk på gatan på en kvartersfest.
Två flickor är blöta och bakom dem står en kvinna som håller ett öppet paraply.
En kvinna i vitt håller i en bukett rosor.
En ung kvinna i "street kläder" och stövlar vid en sjö som utför en balett drag.
En man och en kvinna går uppför en stentrappa och tittar på en videokamera.
Fyra män klädda i t-shirts och shorts tittar ut genom ett fönster till gatan nedanför.
Flera män som står på en parad flyter genom en gata full av människor.
En rynkad gammal man med vitt hår sitter framför ett kedjebundet stängsel.
Skjortlös man skateboard gör trick på en skatepark.
En man med hörlurar går förbi en vägg med röd och lila graffiti.
Två män som bär sombrero's i New York City.
En dam i lila topp och en vit kjol tittar på en marscherande parad.
En person rider en motorcykel nerför en gruskulle.
En kvinna i gult med en barnvagn, och en man i en blå skjorta med en ryggsäck går på en upptagen stad kvarter.
En man i sitt vardagsrum funderar på att packa för en resa.
En afroamerikansk kvinna sitter vid ett brunt bord, klädd i lila klänning, rosa skor och svarta solglasögon.
En man smög in i en stol på en strandpromenad.
Två män, en man som säljer frukt, den andra inspekterar frukten och samtalar med säljaren.
En man och en kvinna kramar på en gata.
Många människor på en stadion klädd i vitt samtalar med varandra.
Många människor har samlats för att titta på något som inte finns på bilden.
Ett par sitter på en bänk och pratar, medan en kvinna går med en hund i bakgrunden.
Två kvinnor i fläckiga klänningar som går på en trottoar.
En grupp flickor leker i en vattenfontän i solen.
Folk landskapsarkitekter och trädgårdar runt gångvägen.
En flintskallig man i röda solglasögon klädd i en grön skjorta som står framför en byggnad.
En barfota pojke med en blå och vit randig handduk står på stranden.
Ett par och två flickor tittar över ett tydligt räcke.
Människor i en produktionsbutik plockar produkter att köpa
En tatueringskonstnär som använder tatueringsfärg på huden.
En kvinna som står bredvid två personer pekar mot himlen.
Ett par går nerför en ö i en butik och säljer konst- och historieböcker.
En man med namnbricka sitter i en stol.
En man på avstånd av ett buddhistiskt tempel.
En man balanserar en metallkula på armen.
En negerhane i vit t-shirt och en svart hatt som sitter på trottoarkanten och sms:ar.
En pojke i svart skjorta bär en blå hink medan han går med män klädda i vitt.
En ung mörkhårig kvinna med rött solskydd som håller ett öppet vitt paraply mitt i en folkmassa
En man som håller i ett litet barn som bär ryggsäck.
En ung man sätter upp biljardbollar, på en lila filt biljard.
Flickor sitter med händerna på knäna
En flicka i en svart tank med shorts till vad som verkar dansa med flera människor runt.
En pojke och flicka i svarta overaller står vänd mot en flicka i rosa jacka, med vuxna i bakgrunden.
En man och en kvinna som knuffar barnvagnar går förbi några människor som säljer föremål i tält.
En kvinna i randiga strumpbyxor vägleds med strängar.
En byggnadsarbetare i en orange väst lägger kullerstenar.
En asiatisk kvinna som sitter utanför ett marknadsstånd.
En man sitter på sitt rum utan att äta i flera dagar.
En husvagn kör ner för en röd tegelväg.
En ung kvinna med brunt hår och tanktopp tar en bild med en kamera.
En person som ligger på en bänk framför en vattenfunktion.
En leende ung man som går på bredvid stranden med baseballmössa, blå t-shirt och jeans.
En grupp människor vinkar till en person på en balkong.
En uniformerad man i armén utbildar en schäfer med armskydd.
Ett barn på skridskor ramp övar coola rörelser.
Vissa män verkar diskutera något på en båt eller ett skepp.
En man med flygmössa och glasögon sitter på vägen.
Folk korsar en trädkantad gata framför en byggnad.
En man i grå skjorta vilar huvudet på ett bord.
En man i vit skjorta och mörka shorts arbetar utomhus.
En kvinna i svarta byxor tittar på sin mobil.
En ung kvinna i rosa skjorta som försöker repa en kalv på rodeon.
En familj står utomhus en molnig dag.
Ett mycket litet barn sitter i handfatet med färg på kroppen och ansiktet och leker med köksblandaren.
Barn som snurrar runt i en glasspinner.
En man och en kvinna håller upp skyltar vid en protest.
En kvinna som jobbar på däck i helgen.
En äldre man, som bär marinblått, sitter på en bänk längs gatan.
En kvinna tar en bild med sin kamera.
En äldre man i blå jeans och brun rock vilar mot en orange byggnad.
En man, hand på huvud, betraktar en Bank of America reklam.
Två kvinnor sitter på en bänk på natten framför en butik
En man i vit skjorta sitter på en låda.
En äldre man med tatueringar och biker regalia dröjer ett ögonblick på en stad gata.
En man sitter ensam och fiskar längs strandlinjen.
En äldre man sitter utanför på en bänk framför en stor banderoll som säger: "Memoria Justicia Sin Olvido."
En man på en cykel i grå jacka bär bladverk.
En pojke med glasögon med en ljusgul skjorta står på en parkeringsplats.
Två män går längs en grusväg.
En mor i blå bast och blå skor med sina två söner.
Två hundar leker med en blå och grön boll.
En man som bär en ljus, flerfärgad hjälm sitter på en motorcykel.
En man hukar sig framför en gul vägg.
Ser ut som en bondemarknad, några tabeller med olika objekt visas.
En blond pojke i blå skjorta sitter med en kvinna i glasögon.
En man i en elegant vit skjorta blickar in i kvinnans ögon medan hon håller i sig på baksidan av sin svarta och rosa klänning.
Folk leker i en fontän vid skymningen.
Fyra pojkar poserar medan en pojke sätter ner sin drink.
På en livlig gata bär en dam gods på huvudet.
En gatuartist i en orange overall rider en lång enhjuling som en publik klockor
En person som sitter på stolen framför en folkmassa.
En hane väntar på att tåget ska anlända till perrongen.
Tre vita män i t-shirt hoppar upp i luften.
En sångare som gör en scendykning i publiken.
En dykkurs som tar en bild under lektionstiden.
En kvinna i randig skjorta viker armarna medan hon står i en livsmedelsbutik.
En trasig bil med många brandmän som skär in i bilen.
Flera människor väntar på att checka ut i en butik med ett lager ser tak.
Två tjejer spelar volleyboll, en slår bollen.
En äldre man häller upp något ur en påse i vattnet.
Sex personer är i en gymnastiksal och arbetar på att reparera några cyklar.
Två unga asiatiska pojkar sparrar med varandra.
En kvinna förbereder ingredienser för en skål soppa.
Två män med shorts jobbar på en blå cykel.
En man och en kvinna som tar en tupplur på en tillfällig rip.
Det finns en man inlindad i en filt av något slag som glider nerför en kulle som är täckt av snö.
En man och kvinna njuter av middag på en fest.
En nationell vaktsoldat leder en grupp andra nationella vaktsoldater som sjunger nationalsången.
Två ungdomar går nerför en lutande gata.
En kvinna på en restaurang dricker ur en kokosnöt och använder ett sugrör.
En kvinna med blå uniform står och tittar ner.
En man i shorts pratar med en annan man i blå jeans framför ett handfat.
En man som matar ett barn i en barnstol.
En ung hjälmcyklist i blått tar upp i luften medan han går över små kullar.
En liten bebis i rosa hatt som ligger naken och sover.
Två barn på magen låg på marken under en pipa.
Två personer pratar i närheten av en röd telefonkiosk medan byggnadsarbetare vilar i närheten.
En infödd kvinna arbetar på ett hantverksprojekt.
Barn jagar bollen i en fotbollsmatch.
Två barn hoppar på en screenad i blå och svart studsmatta medan utanför omgiven av träd.
Två hundar springer på ett fält och tittar på en osynlig frisbee.
En trummis och gitarrist spelar en show i ett mörkt område.
En trio av människor vandrar genom en mycket snöig stig.
En grupp människor är nära en liten flod mitt i en stad.
En kvinna kikar in i ett teleskop i skogen.
En liten blond tjej med en prickig tröja ger ett uppstoppat djur ett "bad" i ett handfat.
En ung man med näsring borstar tänderna.
En snöåkare flyger genom luften, medan andra skidåkare går uppför bogseringsrepet och tittar på.
Tre flickor rider med fokus på den yngsta flickan.
Heavyset kvinna blåser sitt hår med en hårtork leende alla glada
En kock som arbetar i ett kök med kniv.
En man som rör på sig blommor medan en kvinna ger honom en gest.
En kvinna som sjunger i en mikrofon medan en man spelar trummor i bakgrunden.
Mannen som bär mössan ger en nyfångad fisk till pojken i den lila hatten.
En arbetare som klänger sig fast vid ett träd.
Flera människor står runt en skål, där en man manipulerar ett brunt föremål.
En rullskridskomunk med några fina solglasögon ber innan han gör några sjuka tricks.
En kvinna som bär solglasögon och en blå skjorta, som säljer snäckskal, ser på en äldre man med svart skjorta och mössa.
En gammal man sopar golvet när en dam går bort från kameran.
En man med dreadlocks leker med håret på en kvinna som sitter på en stol på en kullerstensgata.
En man arbetar på en byggarbetsplats.
En man är mitt uppe i en röd, vit och blå volleyboll.
En man står i ett rörligt matstånd och tittar ut genom halvdörren.
En basebollspelare med en röd hjälm och vita byxor är taggad av catcher medan du springer till hemmabas.
En man i orange rock sveper ut.
En man i lila skjorta som jobbar i ett biologilabb.
En man leder två små ponnyer på en promenad i en park.
2 kvinnor, 1 från Tyskland och 1 från Kina, tävlar i en brottningsmatch på en matta.
En man och en kvinna som sover på en bänk.
En man och en kvinna sitter på golvet framför bagaget.
Enrickshaw-operatör väntar på sin nästa kund.
Två flickor sitter vid ett bord och arbetar med pysselprojekt.
En man springer genom snön med hjälp av snöskor.
En dansare i röd kostym hoppar upp i luften.
En man är parkerad i en renhållningsbil.
En skäggig man i en tung jacka sitter i ett hörn med en pappersmugg.
Man på en skateboard, med en tom pool som ramp på en mycket vacker dag.
En man med en stor hatt i buskarna.
En närbild av ett barns ansikte som äter en blå hjärtformad klubba.
En man och en kvinna jobbar på att byta ut ett cykeldäcksrör.
En ung pojke visar sitt bruna och gröna pärlhalsband.
En man i grå t-shirt arbetar bälgen för att starta en eld på en tegelugn inuti ett träskjul.
En kvinna som står framför träd och ler.
Någon i asiatisk kostym sitter ner och håller ett svärd.
En ung fotbollsspelare ställer upp för ett field goal.
En kille i en ljusgrön huvtröja går över en korsning medan han tittar på en olycka mellan några bilar och en cykel.
En ung man gör sig redo att sparka en fotboll.
En tävlingslöpare som tar sin första sprint i en tävling.
Två män, en i blått och en i rött, tävlar i en boxningsmatch.
En grupp vänner låg utspritt på golvet och njöt av sin tid tillsammans.
En stående man håller en mikrofon framför en man som håller i en gitarr.
Roller derby flicka skridskor med andra.
En kvinna som hämtar en påse i en affär.
Två motorcyklister tävlar om nacke och nacke runt ett hörn.
En man som står ensam på trottoaren och justerar hatten.
En man med funktionsnedsättning som inte har ben går med en annan man som går in i ett maraton.
Flera kroppar kolliderar i en fotbollsmatch.
Två personer, en klädd som en nunna och den andra i en roger smed t-shirt, kör i en fot ras förbi åskådare i ett skogsområde.
Tre män på hästar under ett lopp.
En mörkhyad man i vita skjortor och en svart ärmlös skjorta kastar sin skateboard på en cementyta omgiven av höga byggnader och palmer.
En man, klädd i en tröja med huva, sitter vid en fontän och tittar på folket i staden.
Simmare står på olika nivåer i ett stort dykbordskomplex i ett rum med figurer från mytologi målade på väggen.
En ung indianpojke som sitter ner och tänker på sin framtid.
En pojke i en huvtröja kastar ett föremål i en smutsig simbassäng.
Färgglada kostymerade män i en föreställning.
Två boxare är redo för sin kamp när publiken tittar med förväntan.
Barn spelar en sport på en plan.
En kvinnlig artist sjunger och spelar gitarr framför en mikrofon.
Pojkar tävlar i kampsporter.
En grupp svarta som uppträder i orangea skjortor framför en inhägnad park.
Skolflickor i uniform marscherar i en parad medan de spelar flöjtliknande instrument.
En man stoppar en fågel från ingredienser i en blå skål.
Pojken hoppar i sin säng med en karatespark.
Ett barn i en hoppstol och en stående pojke omgiven av leksaker.
Det är folk som samlas runt bordet och spelar Jenga.
Jag ser en skäggig man och en äldre dam dela en skål med mat.
En ung man åker skateboard på en cementvägg.
Människor som seglar på en sjö med solen genom molnen i fjärran.
Två män som bär kampsportkläder utövar kampsport.
Ett pojkband och ingen matchar någon borde ha skickat ett PM.
En grupp go-cart ryttare tävlar runt en go-cart spår.
En person klädd i vinterkläder poserar med en snögubbe omgiven av snötäckta landskap.
En man håller en presentation framför en publik.
En medelålders man tejpar knät på en yngre fotbollsspelare som sitter på ett träningsbord.
En tatuerad man i overall på en scen som håller i en mikrofon.
En liten flicka leker med en liten elektrisk krets bestående av tre glödlampor och ett batteri.
Mannen som bär blå hjälm smälter samman med trafiken på en cykel.
Ett gäng unga vuxna stirrar i koncentration på sina datormonitorer när de tävlar.
En ung pojke i gröna övningar jonglerar på en parkeringsplats.
En liten flicka i en prickig klänning ser tillbaka på en kvinna i svart klänning.
En man justerar motorn på en båt nära vattnet.
Det är en tennismatch som spelas på natten i denna stadion.
En barn snowboardåkare kommer till ett stopp
En fotbollsmatch spelas som två män försöker nå bollen innan deras respekterade motståndare.
Unga kvinnor och barn i en by, med en ensamstående kvinna fokuserad på kameran.
Toddler i en grön skjorta borstar tänderna med en gul tandborste, medan mamma övervakar honom.
En man i rullstol och bär en röd joggingdräkt bär en fackla.
En son och hans föräldrar tar en gruppbild i en kyrka.
Tre män tävlar i ett hinderlopp.
Två män observerar en annan när han lägger sista handen på våt cement.
En soldat tittar på kikare i det bergiga landskapet.
En grupp unga pojkar tävlar en snöig dag.
En man hoppar rep medan en massa människor tittar på honom.
En ung pojke och flicka skrattar tillsammans när flickan håller upp en hand skylt.
Två män i motståndarlag tävlar mot en fotboll.
En cyklist som bär en gul skjorta drar av ett otroligt trick i luften.
Två kvinnliga kickboxare, en med lila sportbehå, slåss ut på en arena.
Två män på snabb motorcykel kör runt ett hörn på en kapplöpningsbana.
Två män vaktar mannen med basket under en match i skymningen.
En man som bär ridkängor och hjälm rider en vit häst, och hästen hoppar ett hinder.
En grupp män i kostym spelar musik.
Man och kvinnor tittar genom mjölk lådor fulla av skivor eller bilder på rea.
En tävlingskatamaran lyfts upp på ett skrov i vattnet.
En grupp marinsoldater går längs vägen med amerikanska flaggor och andra militära flaggor.
En man som håller ett dricksglas i kameran.
En man på scenen, spelar gitarr med ljus i bakgrunden.
Fyra unga barn leker med tomma behållare.
En grupp arbetare lyssnar på instruktioner från en kollega.
En tempelridare rider en stor grön traktor nerför vägen under en parad.
Tre hundar leker i vattnet.
En man spelar en trumma och en liten pojke träffar sin egen, lilla trumma.
En grupp tjejer som spelar ett spel på hästryggen.
En man som ser på när en kvinna avfyrar ett vapen med ett leende på skjutavstånd.
Cykelledaren trampar för sitt liv när konkurrerande länder vinner hans svans.
Ett lag av fotbollsspelare är hopkokt och har en seriös diskussion.
En grupp människor i lila skjortor och bruna byxor alla går i samma riktning.
En man i en ljus skjorta spelar trumpet.
Killen med jeansshorts är i skateparken och gör tricks på sin cykel.
Mor och dotter bär Alice i underlandet seder poserar för en bild.
En liten pojke som använder en borr för att göra ett hål i en träbit.
Två cyklister tävlar mot varandra på en grusbana.
En frisbee kastas till flickan medan den andra tjejen verkar be om det.
En ortodontist arbetar på en patient, medan en man håller ljuset.
Två personer äter hamburgare på gräsmattan stolar medan en tredje dricker en burk läsk.
Två bicyklister rider nerför gatan förbi folk medan de pratar.
I en bowlinghall håller en man i svart skjorta en bowlingboll och tittar nerför banan.
Två män i svarta kläder med blå och röda bågar uppträder framför en publik.
Två män, en svart och en vit, spelar sina gitarrer och sjunger in i mikrofoner när de står utomhus.
En kickboxare landar ett flygande knä i ansiktet på sin motståndare.
Tre personer tävlar runt ett rött spår.
Fotbollsspelare kämpar för att få pjäser genom en tuff linje.
Flera män ber medan de står vid slutet av ett matbord.
Två indiska barn i formell dräkt som gärna utför en rituell dans.
Tre barn står nära varandra och bredvid en lång blå trästolpe.
En grupp människor springer.
Två kvinnor går nerför stranden och bär brädor och flippers.
En pojke sitter på en klippa och tittar på dalen nedanför.
En kvinna som står på en hög klippa på ett ben och tittar över en flod.
En brunettkvinna står på trottoaren och tittar nerför vägen.
En grupp av tre vänner samtalar inne i ett hem.
Två kineser står vid en kritbräda.
En person som bär blå jeans och en röd tröja vi vänder hörnet av en tegelvägg.
Jordbrukarna utför sitt jordbruk under dagen.
På någon sorts karneval gör en man sockervadd.
Ett gäng poliser står utanför en buss.
En äldre vithårig kvinna tittar i registret och genom sina glasögon.
Två män står i telefonkiosker utanför.
Två kvinnor klädda i rött och en man kommer ut ur en hamn-a-potty.