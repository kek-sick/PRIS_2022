Två unga, vita män är ute i närheten av många buskar.
Flera män i hårda hattar använder ett jättelikt trissasystem.
En liten flicka som klättrar in i ett lekhus i trä.
En man i blå skjorta står på en stege och städar ett fönster.
Två män är vid spisen och lagar mat.
En man i grönt håller i en gitarr medan den andra mannen iakttar sin skjorta.
En man ler mot ett uppstoppat lejon
En trendig tjej som pratar på sin mobil medan hon glider långsamt nerför gatan.
En kvinna med en stor väska går förbi en grind.
Pojkar som dansar på stolpar mitt i natten.
En balettklass på fem flickor som hoppar i sekvens.
Fyra killar tre bär hattar en inte hoppar på toppen av en trappa.
En svart hund och en fläckig hund slåss
En man i neongrön och orange uniform kör på en grön traktor.
Flera kvinnor väntar utanför i en stad.
En dam i svart topp med glasögon strör pulversocker på en bundt kaka.
En liten flicka sitter framför en stor målad regnbåge.
En man lägger sig på bänken där en vit hund också är bunden.
Fem personer sitter i en cirkel med instrument.
Ett gäng äldre kvinnor spelar sina klarinetter tillsammans när de läser av noter.
En stor struktur har gått sönder och ligger på en väg.
En stor skara människor står utanför framför ingången till en tunnelbanestation.
En man som får en tatuering på ryggen.
Två barn sitter på en liten såg i sanden.
En man som bär en reflekterande väst och en hård hatt håller en flagga på vägen
En person klädd i en blå rock står på en livlig trottoar och studerar målning av en gatuscen.
En man i gröna byxor som går längs vägen.
Det lilla barnet klättrar på röda rep på en lekplats.
Du vet att jag ser ut som Justin Bieber.
En ung man i svart och gul jacka stirrar på något och ler.
En man som står vid en urinoar med en kaffekopp.
Fem personer går med en flerfärgad himmel i bakgrunden.
En gammal man som tar en öl ensam.
En utbildad polishund sitter bredvid sin handledare framför polisbilen.
En person som cyklar på en snöig väg.
Fem män, jämnt klädda i vita skjortor, slips och svarta byxor samtalar på baksidan av en öppen van.
En man med baklängeshatt jobbar på maskiner.
En svart kvinna och en vit man som arbetar i en fabrik och packar burkar med ljus i lådor.
En asiatisk man som sopar gångvägen.
En man lutar sig in i en bil för att tala med föraren, som en man på en cykel ser på.
Två små barn ute på gräset.
Folk tittar på en person i en konstig bil i en plaza.
En man går förbi ett silverfordon.
En vacker brud som går på en trottoar med sin nye man.
En liten pojke som spelar GameCube på McDonald's.
En vit hund skakar på kanten av en strand med en orange boll.
En grupp människor som grillar på en park.
En man i solglasögon lägger armen om en kvinna i en svart och vit blus.
En man med ballonghatt och folk som äter utomhus vid picknickbord.
En pojke hoppar sparkar över tre barn sparkar trä under en tae kwon do tävling.
En pojke i röd jacka som häller vatten på en man i vit skjorta
En man med en röd jacka skyddar sig mot solen när han försöker läsa ett papper.
Män som går nerför en gata med barn.
En liten pojke står på gatan medan en man i overall arbetar på en stenmur.
En svart hund hoppar över en stock.
En man i kostym springer förbi två andra män, även klädda i kostym.
En man i röd skjorta som cyklar runt vattnet.
En barfota man som bär olivgröna shorts grillar korvar på en liten propangrill och håller en blå plastkopp.
En hund springer i snön
En publik står och väntar på grönt ljus.
Man på skidor tittar på konstverk till salu i snön
Sju klättrare stiger upp i ett stenigt ansikte medan en annan man står och håller i repet.
Den unga gymnastens smidiga kropp svävar över balansbalken.
En ung pojke knuffar en leksak ATV runt en gummipool
Kvinnan i röd vindjacka ser ut som en kikare på taket i staden nedanför.
En man står framför ett litet rött föremål som ser ut som ett plan.
En hund leker med en slang.
En man och en liten flicka poserar gärna framför sin vagn i en stormarknad.
En vit hund är på väg att fånga en gul hund leksak.
Killen i grön skjorta med handtäckning en del av ansiktet i restaurangbåset.
En svart och vit hund hoppar upp mot en gul leksak.
Två vandrare vilar vid en snöplätt.
En man som visar upp sin nya träskapelse.
En äldre far och hans vuxna son förbereder sig för en campingtur i vilt tillstånd.
En skäggig resenär i röd skjorta som sitter i en bil och läser en karta.
En ung pojke vinkar handen mot ankan i vattnet omgiven av en grön park.
Ett par sitter på gräset med barn och barnvagn.
Några män står framför en byggnad bredvid en parkerad bil.
Den svarta hunden rinner genom vattnet.
En man borrar sig genom den frusna isen i en damm.
Två stora bruna hundar leker längs en sandstrand.
En person i blå och röd is klättring med två picks.
Tre personer går på en stig på en äng.
En man i svarta kläder skyfflar snö in på gatan, utan hänsyn till all allmän säkerhet.
Ett par står bakom sin bröllopstårta.
En våt svart hund bär en grön leksak genom gräset.
Byborna säljer sina grödor på marknaden.
I en fullsatt konsert närmar sig en vit man huvudsångaren som bär en gul skjorta.
En pojke hoppar på sin skateboard medan en publik tittar
En man och en bebis är i en gul kajak på vatten.
Två personer sitter på en bänk och en kvinna står vid deras sida.
En byggarbetsplats på en gata med tre män som arbetar.
Två män sitter på en bänk och pratar, med en reklamskylt för glasögon i bakgrunden.
En grupp ungdomar marscherar längs gatan och viftar med flaggor som visar färgspektrat.
Tre gamla män ser på när en annan man lagar fisk.
En kvinna i en vit tank topp med en grön strömmande kjol, på scenen sjunga en sång.
Två män och två kvinnor sitter på trappan utomhus.
Ett brunt och svart labb är ute och det svarta labbet fångar en leksak i munnen.
Hockey målvakt pojke i röd jacka hukar efter mål, med pinne.
Mannen med ryggsäcken sitter på en gårdsplan framför en skulpturläsning.
Toddler i en röd hatt som håller i några räcken.
Tre hundar står på ett gräsfält medan en person knäböjer i närheten.
En man står framför en skyskrapa
En kvinna går sin baby med en barnvagn i den lokala parken.
En man i röd skjorta sitter vid frukt till salu.
En ung blondhårig pojke och en mörkhårig flicka äter vid ett barns bord.
Pojken äter sin mat utanför vid bordet.
En svartklädd man spelar elgitarr på en konsert.
En tjej som spelar softball träffar bollen nästan direkt nedåt
En man i svart skjorta spelar en svartfärgad gitarr.
En man som bär en svart skjorta som slätar ut betong i ett stadsområde.
En kvinna i vit skjorta sitter vid ett bord i en trevlig restaurang.
En kvinna ligger på en röd filt i en park.
En ensam man står på en bro på kvällen.
Ett barn går på en gräsbevuxen åker.
En man och hans hund grillar gröna bönor på en grill.
Tre personer vilar på en avsats ovanför moutainerna.
Många människor korsar en mycket lång gångbro med en trädtäckt kulle i bakgrunden.
En ung pojke med utsikt över en skara uppblåsbara båtar.
Två små flickor och en gammal man har ett samtal.
Asiatisk man och blond kvinna håller händer utomhus, man i bakgrunden klockor.
En äldre man med grått hår sitter i en stol och spelar ett stort instrument av bambu.
En man i vit skjorta cyklar på en livlig gata.
En man står på en stege och målar tegelstenar
En 30-årig man som leker med sin telefon på ett tunnelbanetåg.
Två kvinnor går i en korsning med en buss i bakgrunden.
En grupp människor äter knuttor.
En kvinna bär en skål med frukt på huvudet nära havet.
En kille klädd i blått i ett hål.
Fyra barn ler när de poserar tillsammans med en cykel som är alldeles för stor för dem.
Två individer, en man och en kvinna, står i ett skogsområde runt ett badkar.
Ett sovande barn är i någons armar och bär en rosa randig outfit
En medlem av en afrikansk stam tittar uppmärksamt på kameran i stamdräkt.
En samurajkrigare i helsvart klänning tar sitt svärd från skidan på en utomhus träningsmatta.
Flera ungdomar sitter på en järnväg ovanför en fullsatt strand.
Fem vandrare, en vänd mot kameran och de andra vända bort från den, går genom en stenig flodbädd.
En säkerhetsvakt står vid en metall, upplyst skulptur.
Två kvinnor, en i grönt och den andra i lila, som tvättar en trottoar.
Två tjejer hukar sig framför några buskar och pratar på sina telefoner.
En ung flicka bär en flerfärgad håller en orange boll i sin högra hand går genom ljusa grönt gräs bakom ett hus
Ett litet barn som leker med en leksak medan det ligger på golvet.
En liten skateboardpojke gör ett trick på sin bräda medan en annan ung skateboardare klockor.
Två barn skrattar i gräset.
En ung kvinna som håller i en flaska och sträcker ut den från en bänk för att skaka en mans hand.
En förare kommunicerar på sin walkie talkie.
En flicka paddlar nerför en stor flod, sett bakifrån.
En flicka med flätor leker i vattnet.
Ett par bär vita tröjor sitter vid ett restaurangbord.
En måltid ligger på ett bord i en restaurang.
Två byggnadsarbetare sätter sig på en stålbalk.
Ett barn som gärna blandar smet i en skål.
Två barn leker med en ballong i lera en solig dag.
En liten flicka som tittar på en broschyr om tågturer
Två kvinnor sitter och pratar och skrattar tillsammans.
Folk joggar tillsammans på en strandpromenad.
Ett litet barn hoppar från ett högt dyk vid poolen.
En ljusfärgad hund springer på stranden.
En man bor i ett vattenfat av trä och äter en frukt.
En man sover på en bänk nära en busshållplats.
En liten flicka i röd skjorta och jeans klättrar upp i ett litet träd medan en annan liten flicka tittar på.
En man som sover i en bil som kör.
En kvinna i röd skjorta ligger under en filt och sover i ett fordon.
En man i ett hemkök vänder en pannkaka extremt högt.
Flera brandmän svarar på ett larm.
Flera brandmän står utanför en byggnad nära sina brandbilar.
En strand med blå och röda båtar, med människor på stranden
Män som bär hattar och skyddsvästar arbetar.
En tidskriftsförsäljare sitter bakom ett mycket färgglatt collage av tidskrifter.
En man i hård hatt bär en blå skjorta och blå jeans overaller.
På bageriet sover den feta gamla bagaren medan hans lärling gnuggar mjölet ur hans ögon och sitter bredvid honom.
En grupp skjortlösa män sitter i skuggan på en tropisk strand.
En pojke i sina blå badbyxor på stranden.
En skidåkare har utsikt över ett snötäckt berg.
En pojke som bär en röd skjorta cyklar bredvid en hög med smuts.
Cyklare i ett cykellopp tar en skarp vänstersväng.
Tre pojkar leker och cyklar med en sandhög i mitten
Äldre man med käpp böjer sig över nära en man och kvinna.
En läkare och sköterskor i blå skrubb utför en operation.
En svart och vit hund hoppar efter en gul leksak.
En ullig hund jagar en doberman på en strand.
En man står där efter att ha rullat en bowlingboll nerför en fil.
En gammal, uttorkad, skäggig man klädd i svart, ridande på en vacker vit åsna på vita klippor.
En man och en kvinna som sover på en blå soffa.
En man i gul skjorta kastar ett spjut på ett spår.
En publik tittar på luftballonger på natten.
En kvinna läser en tidskrift över en annan kvinnas axel.
Två män på huk för att tända ljus på natten.
En ung man går genom en livlig gata vid ett köpcentrum.
Den lille pojken cyklar i ett lopp.
En grupp människor som sitter vid ett bord i ett mörkt rum.
En man med två hundar på en strand
En pojke som är täckt av suds har rengjort ansiktet.
Dussintals människor festar på en båt.
En ung kvinna på en båt i en ljusfärgad bikini sparkar en man i en halmhake.
En pojke glider ner för en bild i en pool med färgglada rör.
En man i våtdräkt kastar upp ett litet barn i luften och är redo att fånga honom.
En grupp människor som rider i baksätet på en lastbil, längs vägen, i ett landsområde.
Två kockar lagar hamburgare i ett restaurangkök.
Två unga pojkar gör löjliga ansikten.
En person med bruna byxor sitter runt ett inhägnat område som har gnistor som flyger.
Kvinna på en kulle vid ett vitt kors med utsikt över en strand.
Fyra flickor sitter i gräset medan flera män står nära dem.
Män på jobbet skyfflar snö från ett järnvägsspår.
En man, en flicka och två hästar är nära en innesluten eld.
Arbetare med reflekterande västar som arbetar nära en tågbil.
En äldre kille tittar på en klassisk, rustik, volkswagen skalbagge.
En kvinna sätter ihop en vit metallram på trottoaren.
Det finns tre hundar som stirrar på en boll mitt i dem.
En skjortlös man och en kvinna som sitter på en docka.
Män i skyddsvästar jobbar på ett spår.
En man som fixar vägen med sin utrustning.
En kvinna med rött hår applicerar mascara på sina ögonfransar.
En vit hund har huvudet på marken.
En kvinna i blå shorts och en vit skjorta är inomhus bergsklättring.
Många skotrar parkeras tillsammans på trottoaren.
Parkens polishelikopter förbereder sig för landning.
En man i en reflekterande jacka ställer sig på ställningen.
En grupp på fjorton personer samlas i en sal med matbord och en scen.
En tonårspojke hoppar på en uppblåsbar bild.
En familj som leker på en traktor en vacker dag
En äldre kvinna steker mat i ett kök.
Två unga människor blir närda av en praktfull ung kvinna klädd i en röd bikini och en röd fjäderklädd huvudbonad.
Två skidåkare tar sig genom skogen.
Skidåkare på toppen av en snötäckt kulle.
En brun hund som springer bredvid gräs.
En kvinna i grön skjorta och jeans knäböjer på en toop med kaffe i handen, hennes handväska bredvid henne och en stor dörr bakom henne, när hon fyller i pappersarbete.
Folk korsar en gatukorsning.
En kvinna klädd i ljuslila och klädd i en korsage knäpper händerna i knät.
En mor och barn fiskar på en strandpromenad på natten.
Sex män spelar ett spel i sanden med träpaddlar.
En kvinna i en grön tanktopp är omgiven av tre barn som skrattar.
En man i svart skjorta, och svarta byxor, arbetar på motorn i en gammal, grön antik bil, med en gul gasbehållare sitter på gräset.
En kvinna i en blå jacka rider en brun ponny nära vattnet.
Två hästar drar en vagn som körs av en kvinna över snötäckt mark.
En person som klättrar nerför en klippa med hjälp av ett rep
Gruppen av vandrare vilar framför ett berg.
En kvinna som står framför en kritritning
Tre unga vuxna sitter här och tjejen låtsas sparka en av killarna i ansiktet medan han skrattar, och killen bakom honom ser ut som om han är mitt i natten.
En grupp barn i klassen med händerna i luften.
En man som bär badbyxor hoppar från en betongplattform ner i en stor vattenförekomst.
Kvinnan arbetar minutiöst med en symaskin.
En dam i vit t-shirt tittar mot personen med armen upp i luften.
En tjej som jobbar på en gårdsmarknad och säljer paprika.
En äldre kvinna sitter i en stol med en käpp i handen.
En pojke har blåst fyra bubblor på gräsmattan.
En liten pojke som leker i vattnet.
Hunden får slut på tunnel på hinderbana
En gul hund och en svart och vit hund springer i smutsen.
Två män barbecue på en strand.
En liten flicka i en blomtrycks baddräkt, hoppar i havet.
Lilla flicka i blå baddräkt står på en ledstång nära en strand.
En ung asiatisk pojke sitter på ett räcke bakom en rad färgglada hattar
En vit och svart hund hoppar in i en pool.
Pojkarna ler under vattnet vid poolen.
Två personer som har en diskussion sitter i en restaurang.
Flera personer tar en paus på en snöskotertur.
Två personer arbetar på att ta bort snö från ett tak.
En ung man i svart skjorta tar en fällstol från en stor hög.
En kvinna går i skymningen nerför en stadsgata.
En liten flicka med brunt hår blåser bort kronbladen från en blomma.
Tre personer på ATV är utanför.
En man på en fyrhjuling flyger genom luften.
En man på en fyrhjuling hoppar nära en liten byggnad.
En kvinna med mörkt hår i bikini sitter på en strand.
Två händer vänder lite mat i en gjutjärnspanna, med en spatel.
Två kvinnor kramas i en gräsbevuxen, inhägnad åker med en ko bakom i bakgrunden.
Ett stort skepp närmar sig hamnen med två män som väntar på dess ankomst.
En man i sandaler och vit kofta sitter på en grön bänk medan han pratar på sin mobiltelefon.
En man på scenen som sjunger in i en mikrofon.
Tre killar rider på en elefant med husliknande strukturer och träd i bakgrunden.
En mexikansk man sitter under motorhuven på sin lastbil.
En pojke i gula glasögon och rödhårig flicka poserar för kameran.
En grupp människor samlas och håller olika typer av flaggor.
En vit pojke som gråter över en spetsig leksak.
En liten pojke bär en fotbollsboll på ett fält.
En kvinna tittar på när en kille tar glass från en frys.
En grupp människor sitter på pallar och äter lite mat
Folk står runt en amerikansk flagga som är utspridd, vänd åt fel håll.
En ung flicka som målar en bild.
En cyklist cyklar på en svängd väg uppför en kulle.
En liten flicka i en jeansjacka som springer genom ett fält.
Mannen i blå skjorta och svarta byxor tittar på tummen på ena handen medan han håller glasögon i den andra handen.
Ett par kysser när de går upp i rulltrappan.
En fotbollsspelare i en grön uniform med en boll i är händer hålls upp av några av sina lagkamrater, medan en motståndare i rött sträcker sig för bollen.
Män bygger en mur i öknen.
En ung grupp vänner prydda med ansiktsfärg och fjäderklädda pannband sitter på en bänk.
Damen har en svart slangväska.
En man i svart jacka står med en grupp människor bakom sig.
En svart hund hoppar för att fånga en rep leksak
En ung flicka tittar genom en gammaldags videokamera.
Flickan i udda kläder läser en broschyr medan hon sitter på en veranda i trä.
En man klädd i en funky outfit spelar gitarr.
En hockey målvakt försöker förhindra ett mål från motståndarlaget.
En vuxen och ett barn går längs stranden under dagen.
En man i förkläde sitter på en trottoarkant.
En brun och vit hund hoppar upp för att fånga en frisbee medan en publik tittar.
Två tennisspelare pratar på tennisbanorna.
Två jonglörer som använder flammande facklor uppträder för en skara människor som sitter på trappan.
Två barn som springer utan skor.
Ett barn sitter på och leker med släta stenar.
En pojke i en Gap-hatt gör ett dumt ansikte.
Fem män, en klädd i en vit skjorta stående på något, hängande upp en bild av ett barn.
En person i hatt leker med en pojke på en strand.
En tjej i en grön Speedo topp och blå goggles håller andan under vattnet.
Pojkar på en motorskoter som rider på en livlig stadsgata.
Två damer och en man som spelar kortspel och dricker öl.
Folk njuter av en samling med Pabst Blue Ribbon och Diet Coke.
Man med röda skor, vit skjorta och grå byxor klättring.
En bergsbestigare klättrar upp för en stor klippa.
En liten flicka som leker i vatten på en grodskulptur.
En hund springer på stranden.
Folk som sitter på en restaurang och äter och man läser tidningen.
En tjej som bär en röd kort och en vit skjorta som tittar genom ett hål.
Svartvit fågel står på handen av någon som håller solrosfrön
En kvinna i vit skjorta och rosa kjol är på väg att träffa en tennisboll.
En hund står i sanden.
Det här är en man som står på ett tak med konstruktion i bakgrunden.
En man tittar genom en stor kameraliknande apparat i ett fält nära en husbil och några parkerade fordon.
En liten pojke står och surfar.
En kvinna i muslimsk klädsel går med en ung pojke längre ner på gatan.
Den lilla hunden springer över gräsmattan.
En kvinna joggar på en trottoar bredvid en högt uppsatt gräsplattform.
En man i röda byxor som hoppar på ett parkbord.
En hund med munnen öppen springer genom ett fält mot kameran.
Smickrande lilla flicka som simmar i utomhuspoolen.
En cykel som sitter på en gata med ett rep bundet till den och en kille som går på repet.
En man och ett barn på ett skepp som sköter underhållet.
Ett litet barn som gör ett handstånd på en säng.
Män med orange skyddsväst arbetar med gatureparationer.
En man med skyddsväst knäböjer och städar tegelstenarna.
Arbetaren håller på att reparera på en gata.
Människan står på vit sand och håller i en snowboard.
En man i orange väst som står ovanpå en byggnad.
En kille i gul skjorta och ljusbruna byxor spelar golf medan publiken tittar på.
En ung flicka i karateuniform med en stor trofé.
Ett barn med flytare som hoppar ner i en sjö.
En kvinna i rosa skär en hamburgare med en spatel.
En pojke i en smutsig skjorta går genom knähögt havsvatten.
En man som står bredvid en naken staty.
Ett litet barn klädd i vitt ler medan en dam hjälper honom att vifta med en flagga.
En person står på en byggnad på sjön.
En ung man i grå jacka står bakom disken i en juvelerarbutik och ler.
Folk går upp och ner för trappan till en kyrka.
Ett antal barn roar sig på kusten av en stad.
En hona jobbar nära havssidan.
Två män arbetar på ett snickeriprojekt med handverktyg.
En kvinna och två flickor klädda i rosa.
En man i svart kostym och portfölj som skyndar sig någonstans, medan han pratar på sin mobil.
En brunettkvinna som går nerför en gata med en kopp.
En skallig liten pojke håller en kyckling medan två män sitter i bakgrunden.
En man som sitter på en vägg och tittar på en vattensamling.
Två hundar springer genom vattnet med ett rep i munnen.
En pojke promenerar vid en damm i en park.
Blond barn med stor svart rock, flerfärgad halsduk, och sticka hatt stående framför ett fönster.
Brun hund med tennisboll i munnen, i vatten och buskar.
Två bruna hundar rinner genom vattnet.
En tjej som blåser bubblor i poolen.
En hög med sjögräs sitter på sanden, bakom den springer en stor svart hund i vattnet.
En ung pojke springer medan han bär sandaler.
En brun och vit hund står utanför medan det snöar.
Någon som arbetar med ett projekt med hjälp av en skärmaskin.
En dams roller derby team tar en paus.
En pojke hoppar från en säng till en annan.
En man i gul skjorta som står mitt i två sängar som en pojke hoppar på i bakgrunden
En ung man med en stor motorsåg.
En man på en motorcykel utan skjorta och en annan man som står under skugga.
Tre personer går in i en byggnad med en handskriven skylt där det står "Välkommen Bikers".
En man sätter upp en mur.
En brunhårig kvinna tittar på ett barn som äter något.
En rad människor, en del stående och en del sittande, väntar på en plattform för ett tåg.
Två skidåkare står, två sitter i backen.
Folk promenerar i ett köpcentrum med färgglada dekorationer hängande från taket.
En kvinnlig smed skor en häst.
Barnet i den gröna kostymen går förbi ett skyltfönster.
En grupp tjejer hejar.
En man är inne i en lastbil och tittar ut med vänster arm framför en dörr.
Ett barn som kliver ur bilen med fotbollsskor.
En vit, ung man i dreadlocks och en grön kilt sitter på en soffa och ler.
En man i blå skjorta kysser en kvinna med blont hår på kinden.
En man och kvinnor poserar för kameran och ser väldigt lyckliga ut tillsammans.
Två barn leker på stigen i en park.
En mycket färgstark buss dras av till sidan av vägen när passagerarna lastar.
En leende kvinna håller en person klädd i en grisdräkt.
En kvinna som bär en blå hjälm cyklar på en parkeringsplats.
En liten flicka i grön klänning står framför pölen.
En man som bär hjälm och cyklar nerför gatan.
Ung pojke och en äldre man som väntar på att få checka ut.
Två personer tar in scenen när de står tillsammans och tittar ut över ravinen.
En kvinna med hjälm som håller i en cykel.
En ung man som står framför en röd godsbil och håller en kamera och tar ett foto.
En person i blå shorts och bär en Walkman joggingspelare.
En man och en kvinna leker på ett träd medan andra ser på.
En grupp ungdomar är i ett garage
Tre män tittar på en skylt på ett kors i en ravin.
En ung dam sitter framför ett stängsel med en hink.
Kvinnan försöker gömma sig under en svart tröja, men hennes röda manchesterbyxor avslöjar henne.
En ung man som städar en staty med en pensel.
Två unga män håller trasor i sina händer, när en äldre man talar om för dem hur de skall rena det stora korset.
En kvinna sitter på en mans axlar med en tung pensel som hammare.
Gruppering av ett träkors nära ett stort stenblock.
En ung pojke plockar upp en pensel och flinar.
Fyra män i vita skjortor och kepsar sitter runt ett bord.
En pojke som tittar på en hackad stock.
Man med grått hår berättar en historia för en grupp yngre människor på en bänk.
Två personer står på ett fält och håller i några böcker.
En person som gör en skateboard vända bredvid en svart soptunna.
En man som står på en järnvägsbana och tittar genom kikaren vid en flod.
Många människor sitter på marken nära en halmhydda.
Ett barn kanske spelar fotboll i kostym.
Människor på cyklar väntar vid en korsning.
En byggnadsarbetare bygger byggnadsställningar för jobbet.
En liten bebis klädd i grönt och gult med ett hakskrik.
En skjortlös man som leder en häst som drar i en vagn.
En kille som står utanför utan tröja och tittar upp på byggnaden.
Den unga flickan svingar högt över marken på en trevlig sommardag.
En ung man gör ett skateboardtrick från en betongbänk.
Mannen håller nätet för pojken som spelar baseball.
En äldre man hukar sig för att lyfta täcket av grillen bär flera shish kabab grillar.
En man med svart skjorta och glasögon springer längs gatan
Ett fempersoners operationsteam är på väg att utföra en operation på ett sjukhus.
En pojke som står på stranden och håller en blå blek och en grön spade.
En liten flicka snurrar i vågorna i den ljusa solen.
Tre personer sitter ute på små stenar bakom en stor buske, klädda i långa byxor.
En man med en högafflar står nära en hink av grenar mittemot ett lägenhetskomplex.
En groundskeeper har samlat en hink full av pinnar.
Svart och vit hund tittar på kameran med mannen böjd över i bakgrunden.
En man som bär hängslen när han står på ett tåg.
Två män och två kvinnor lagar en stor måltid i köket.
Tjejen lär sig om djur på zoo.
En grupp vänner fiskar utanför lastrampen
En mor och son läste en bok om dinosaurier tillsammans.
Två kvinnor, som sitter vid ett bord, med ett grönt sugrör inuti en drink.
En liten pojke i overall som gråter.
Tre män sätter upp en släde på en snöig slätt.
En person sitter bakom två stora brödkorgar.
En man i pilotuniform går nerför trottoaren och bär bagage.
Människor som går längs en flod nära ett vackert hus.
En kvinnlig simmare som bär en badmössa och näsklipp rör sig långsamt genom vattnet syns underifrån.
Fyra män sitter och jobbar på bärbara datorer.
En man i en basebollmössa rensar ut en blåfärgad grop utanför där färgglada julljus hänger ovanför honom.
En flicka som sover med en docka i en prinsessdräkt
En hona tvättar sin medelstora hund utomhus i en plastbehållare medan en vän säkrar den med koppel.
Ett barn som hoppar ner i en vattenpöl.
Barn i svart jacka, röda byxor och fleece hade sovplatser på en röd jacka.
Gubben i brun hatt sitter på bänken.
Tre barn på en gräsplan, en av dem letar efter mat i sin mammas handväska.
En svart man driver en orange trana.
Tre flickor går under en argor på en stig omgiven av träd.
En strand är full av många människor.
Människor samlas runt och promenader köpa en uppvisning av kläder och andra föremål.
Man paddlar en båt på en flod nära stranden.
Två kvinnor står tillsammans och håller i en gryta och en kastrull mat.
En ung flicka med gula flip-flops sitter på ett stort stenblock.
Blond kvinna kör en röd cykel vagn håller toppen av sin hatt och poserar för kameran med en kund sitter i ryggen.
En ung pojke i ett blommigt förkläde hjälper sin mor att laga mat.
En ung man presenterar en annan kvinna med en tårta med tre ljus ovanpå.
Kvinnan med hatten säljer lite frukt och rotfrukter.
Person med en huva jacka sittande på snö framför ett gult tält.
Två hundar brottas på ett gräsfält.
En man i skyddsväst knäböjer och jobbar på ett tåg.
Fem byggnadsarbetare gräver ett hål för att plantera ett träd.
En man i röd skjorta ger leksaker till en liten hund.
Gammal dam som sitter i ett rum fullt av blommor.
5 idrottare bär vita toppar och vita bottnar gör en rutin för en publik.
Byggarbetare står utanför och tittar på ledningar ovanför dem.
En lycklig ung pojke sitter i en stol med en stor Elmodocka.
Ett barn borstar ett spädbarns hår.
Ung man som visar upp sig genom att utföra ett karatedrag för överraskad flicka.
En man som äter i ett stökigt kök.
En tonårspojke har en silverring som sticker ut från näsan.
Den här mannen ler väldigt stort vid kameran.
En grupp ungdomar leker i en källa med vatten.
En kvinna som kastar en frisbee på en strand.
Den mörkbruna hunden leker med den ljusbruna hunden.
En kille som har skyddsutrustning svetsar en stålbalk.
Man i orange shorts bygger ett sandslott, som kombinerar flera bilder till en som resulterar i fyra exemplar av honom.
Två män och en hund står bland böljande gröna kullar.
En grupp människor som går på en gata framför en AMC-byggnad.
En vit man med glasögon blåser en bubbla i ett hus.
En vuxen visar ett litet barn en fäktningsdräkt som sätts upp på ett träd.
En stor hund fångar en boll på näsan
En man och två kvinnor bär alla svarta agera ut en scen framför en byggnad med trappsteg.
Två barn som bär jeans sprutar vatten på varandra.
En brunfärgad hund hoppar in i en utomhuspool.
Folk som sitter i en cirkel med en bok i mitten.
Par, man och kvinna, med liten flicka alla klädda i bröllopskläder medan står längs strandlinjen.
Massor av människor som går under en markis av rosa och vita ballonger
En linje på sex barn i baddräkt förbereder sig för att hoppa in i en simbassäng.
Två bagerianställda som bär röda förkläden håller på att laga mat.
Ett litet barn med röd mössa och en anka är i gräset.
Föräldrar knuffar små barn i röda bilar.
En man i blå skjorta använder en vattningsslang och en annan man i brun skjorta rör på sig presenningar.
Tre pojkar i Florida Marlins hattar.
En familj kommer tillbaka från shopping och en gentlemän läser hans tidning till sidan av gatan.
Två kvinnor som håller händerna i luften medan de hoppar.
En kvinna bär ett barn i armen och håller ett annat barns hand när de går ut bredvid en byggnad.
En hund går genom ett fält.
En livlig gata med massor av människor som står och pratar och två håller i cyklar.
En färgad kvinna som rullar en bowlingboll i en gränd.
En fotbollsspelare i en röd uniform följer efter bollen och kämpar mot en spelare i vitt.
En grupp människor går nerför en stig i skogen.
Tre barn leker med en röd boll i en park.
En liten pojke som sparkar en gummiboll.
Den här bilden av en man som läser är lutad.
En man på en stege klädd i blå jacka och blå jeans
Tre vägarbetare i orangea jackor och byxor städar upp med en skottkärra.
En man på styltor står framför en rad trummisar.
En ung kille, förmodligen i tjugoårsåldern, visar upp sina kulinariska färdigheter med stolthet.
Terrier hund leker med leksak på filt
En hund springer över ett gräsfält med en käpp i munnen.
En pojke med glasögon och rutig skjorta läser en bok.
En ung man tittar på en bok på marken i ett skogsområde.
Två män står i kö på en restaurang.
Flera barn sitter på en karnevaltur framför ansiktet på en clown och flera falska ballonger.
En kvinna med smutsigt blont hår och glasögon skär något.
En man som bär bollmössa och en blå T-shirt rider en vit häst nerför en grusväg genom frodig, grön natur.
En medelålders kvinna som lagar mat medan hennes hund tittar på.
Rödhårig kvinna i flätor och glasögon sy på en symaskin.
Två män i ett rum tittar på en datorskärm.
En grå hund springer längs sidan en pool medan en gul hund hoppar in i poolen.
Ett barn glider nerför en kulle på en släde.
En man och en kvinna som låser armarna (med dyra kläder) bredvid glasdisplayen (kanske butiker) på trottoaren i en urban miljö.
Två arbetare sliter i en smältfabrik.
En gammal kvinna sitter på en transitstation bredvid en bakgrundsbelyst annons.
Folk väntar utanför en byggnad bredvid en väggmålning.
Tre personer knuffar en stor maskin genom gatan.
En man med ärmlös skjorta och bygghjälm.
En man med skägg och hatt tigger pengar från folk.
Flickan på enhjulingen sträcker sig efter barnet på skotern.
Skidåkare åker fast på dammiga sluttningar och faller nästan ner och bryter benen.
En man som bär en plastlapp med en krabba på, håller upp en trähammare.
En man hoppar från en liten stenbro medan tre barn och en kvinna vaktar honom.
Person som sitter på betonglandning bredvid vattenförekomsten
En man som spelar gitarr medan ett par lyssnar och ser en annan man dansa till musiken.
Vissa byggnadsarbetare tar en paus.
En kvinna i en klargrön tröja leker med en drakdocka en trädgård.
Stora mängder människor sitter upp mot väggarna i byggnader.
Ett barn håller gröna skor går i sanden vid vattnet.
En bröllopsdag med bruden i en ljus vit vacker klänning
En person som bär lila jacka står bakom ett högt träd.
Kunderna väntar på service vid en takeout fönster.
En kvinna med blommig skjorta och handväska och en man med svart skjorta går medan en annan man går bakom dem.
Fågelns syn på en man som stiger uppför en trappa utomhus.
Män och kvinnor med vita badmössor som ger varandra turer.
En familj sitter utanför och roar sig i ett parkområde.
En brunettkvinna sitter i en blå fällstol och läser på stranden.
Kommunister rusar för att komma på det sena tåget.
Ett barn och ett litet barn sitter tillsammans i en barnstol.
En grupp tillbedjare håller sina gudstjänster i en offentlig park.
En man sitter framför en datormonitor och håller ett tangentbord och tittar på kameran.
Ett barn ligger ner på en träbänk.
Omgiven av åskådare, en man i röd skjorta, vita byxor och visir, svänger en golfklubba.
Två män diskuterar någon gång nära en vägg med lite graffiti på den.
Vissa personer med svarta bälten, eller svarta och röda bälten, utför kampsporter på en grön matta.
En kvinnlig kampsport student demonstrerar med ett vapen medan andra tittar.
Flera unga vuxna uppträder i kampsportkläder.
En ung kvinna sitter på ett varuhus märkt glass och program.
En pojke poserar för en bild och i bakgrunden hänger en man i ett rep.
Två personer sitter med ryggen vänd mot sockervadd.
En flicka i gul klänning med solen skiner i ansiktet
Åtta herrar arbetar med sten &amp; kakel.
2 kvinnor med färgglada kläder sitter bredvid en grusväg på en sten med en konversation medan de tittar på fältet.
Två män i svart äter en smörgås.
Närbild av en man i en bar, håller sina glasögon lutade framför hans ansikte.
En pojke sitter på rektangulära block.
Ett barn leker på gatan, kör ett hjul.
En man sitter bakom en hård trädisk.
En man i svart jacka tar ett foto på en man i röd jacka.
En man i gul overall ro en båt med en fågel framför sig.
En hane med hatt jonglerar med fyra bollar.
En person i svart hatt håller i flerfärgade jongleringsnålar.
Fem personer sitter runt ett bord, utanför, och spelar ett kortspel.
Familjen sitter på en bänk nära stranden.
En man och en kvinna kan laga mat på lägret tillsammans.
De fyra vandrare gick uppför grusvägen.
Två afroamerikaner gör sina trumpeter i en stor stad med åskådare som tittar.
Folk på avstånd försöker klättra uppför en klippa.
Två poliser tittar på ett hus på avstånd med kikare.
En grupp barn i bruna kläder uppträder.
Två unga manliga vandrare använder en karta och kompass för att hitta sin riktning i skogen.
Två män på en pråm
Tre barn, baby i mitten, sitter i en utomhus swing stol.
Ett barn står redo med en baseballhandske.
Två flickor som står på gräs möter varandra.
Grupp av människor som går på den tunga snön.
Två arbetare som arbetar på sidan av en gata i neongula västar.
Stadsarbetare som sätter betong på en väg.
En byggnadsarbetare som arbetar på flera ställen på vägen.
En man med rött hår som jobbar på sin cykel.
En kvinna som sitter på en bänk framför en stor målning.
En ung pojke spelar på en gunga.
Två män i skogen använder en motorsåg för att hugga några träd.
Byggarbetare arbetar på en väg in i natten.
En man i svart jacka spelar gitarr.
Grupp av människor som står eller sitter utanför ett café.
En man med gitarr sitter på en bänk utanför med tre andra människor som sitter bredvid honom.
En man och en kvinna fiskar från en båt.
Ett litet barn håller en sked i munnen medan det sitter i en stol.
En man i en solbränd fiskares mössa sätter läppbalsam på en kvinna i en båt.
En man justerar rattarna på en stor ljudblandningstavla.
En kvinna i randig skjorta och svart hår står mot några bås.
En svart hund och en brun hund som leker i långa ogräs.
En man i en röd och vit kontrollerad skjorta spelar i en park.
Två män mäter en vägg på en öppen byggarbetsplats.
En man i vit skjorta spelar tennis.
En brun hund som hoppar i luften på en brun slätt.
En ung kvinna som står på en fönsterkant av tegelbyggnad medan barnet tittar på.
Två tonårstjejer, den ena klädd i vit tröja och den andra klädd i röd tröja, spelar fotboll.
En ung bebis som suger en Binky som sover i en stol.
En man som drar en tjusig rickshaw längs en vattenväg ler och ger "tummarna upp" skylten.
En närbild av ett barn på en lekplats med vuxen handledning.
En man i röd skjorta fäster en yngre man i vit skjorta till en blå vadderad matta.
Dessa män utövar kampsport.
Kvinnor och män i ett annat land ser ut som de klappar
En kvinna handlar på en bondemarknad.
Människor går runt och minglar i ett stort öppet utrymme med en hund.
Två kvinnor som bär hattar täckta av blommor poserar.
Den lilla flickan rider i en brun häst.
En tonårspojke pratar med en grupp tonårsflickor.
En man sitter på en utebar nära många läsk och ölburkar.
Tre personer står utanför runt två grillar där kött tillagas.
En asiatisk familj är picknick på stranden medan andra leker i vattnet.
Två män i höga hattar rynkar på kameran
Tre personer sitter på träbänkar på vit och orange kakel.
Mannen bär en vit skjorta och solglasögon.
En grupp på tre personer arbetar i en belamrad kontorsmiljö.
En pojke i våtdräkt hoppar in i en pool med en skallig man.
En pojke dyker ner från en dykbräda i en simbassäng.
Två räddningspersonal är på platsen för en incident.
En man som skapar ett lerföremål vid ett krukmakarhjul.
Folk som grillar vid stranden.
En kvinna håller en liten flicka som försöker fånga bubblor.
Två män hänger och grillar.
En kvinna som spelar gitarr inför en grupp människor som står utanför.
Två hundar leker tillsammans på grönt gräs.
En konstnär konsulterar planen för sin del av en utstuderad kritritning på en trottoar.
En man på jobbet, slaktar en ko.
En man med en stor fjäder i hatten rider en häst.
Två personer bär en stor, uppblåsbar flaska, förbi en ung kvinna och en parkerad vit bil.
Dessa flickor är i uniformer och spelar fälthockey.
En vit och solbränd hund hoppar genom luften.
En kvinna som kastade en bowlingboll i en bowlinghall.
En man spelar trummor medan en annan sjunger Karaoke.
En brun häst står nära en svart häst som sitter på marken.
Ett barn tittar över en karneval monter disk på de olika leksaker.
En man sover i en hängmatta bredvid vatten och en båt.
Elva små flickor poserar som ett lag i en pool.
En man i grå och svart tröja sitter på en pall framför en grupp burar.
En ovanligt klädd man som sitter bredvid en glasskylare.
En man i brun skjorta sitter på trottoaren och spelar gitarr.
En liten flicka med en tiara som äter i någons knä.
En svart och brun hund ligger på en vit matta.
De tre flickorna satt på stranden.
En liten pojke tittar på sin spegelbild i en graverad marmorvägg.
Män och kvinnor på cyklar stannar för att titta på något.
En liten flicka i rosa danser med händerna på höfterna.
En man och kvinna njuter av en cigarett utanför en affär.
En asiatisk stad på natten med ett stort antal människor som går runt.
En kvinna med en blå jacka som sträcker sig ut till ett barn.
En man klädd som kock njuter av en måltid och en flaska vin i en tom restaurang.
En man med ansiktshår i vita kläder som äter en biff.
Tre män arbetar snabbt med att laga mat i köket på en förstklassig kinesisk restaurang.
En man sitter på en sten.
En ung flicka i en gul dans, dansar på en scen med ett basebollfält i bakgrunden.
Barnen leker i skogsområdet nära vattnet.
En flicka i rosa skjorta ligger på ryggen i gräset.
Ett par har ett tecken som visar att de undervisar barn om fred.
Tre personer bär färgglada kostymer och masker som sitter mellan två stenstatyer.
En man på cykel rider nerför en stenig kulle.
Tre unga flickor dansar på stranden i sanden.
Ung flicka i blå klänning kliver över en fotbollsboll.
En snårande brun och svart hund hörn en brun långhårig katt under en trä bänk.
Många människor står och tittar på något.
2 personer sitter barfota i ett tält, en med en öl och en lounging spelar gitarr.
En man i shorts hugger ved utanför en teepee.
En pojke i randig skjorta och en flicka i grön skjorta varje ridning på cyklar med träningshjul.
En vuxen och ett barn sitter på en polis motorcykel.
En man utan skjorta och hatt använder hammare och städ.
En kvinna i svart spelar ett Cello-instrument.
Två män i en träbåt, en klädd i gult och en klädd i svart, färdas på en slät vattenförekomst.
En ung man med ingefära timme spelar en omgång pool.
En man i röd dräkt rider en röd motorcykel uppför en motocross krets.
En kvinna som ger en blondhårig bebis en drink från en kopp.
Sex kvinnor sitter vid ett bord tillsammans framför en bokhylla.
Folk går förbi en uppvisning av underkläder hängande i ett bås.
Två bicyklister poserar av en bäck för en bild.
Två barn står på ett grönt metallstängsel.
En ung pojke med en smart svart och vit skjorta med huvudet böjt
En lastbil har just kraschat i baksätet på en annan lastbil.
Två restauranganställda byter en tallrik mat under en mongolisk BBQ neonskylt.
Två pojkar som leker i vattnet med shorts.
En grön John Deere traktor i ett fält som drar en röd trailer.
Två barn leker på en förskjutningspipa.
En varierad folkmassa kvarnar om (eller grovhus) på en allmän gata, med massor av cyklar på display.
Två personer hoppar jacks på stranden
Det finns ett dussin män i arbetskläder som får vägbeskrivning för en uppgift.
De tre hundarna är på väg nerför gatan.
Damen i den röda bilen går över bron.
En tjej med en svart väska som sitter på en träbänk.
En man i rutig skjorta som kopplar sin svarta laptop till mikroskopet.
En man målar på en trottoar i staden.
En flicka i vit skjorta sitter på en parkbänk med en hund bredvid sig.
En man som cyklar med en grön skjorta med en drink i handen.
En man spelar ett litet gitarrliknande instrument och sjunger in i en mikrofon.
Kvinnorna med shorts har handen på en vit bil.
En person står med ett ben uppstött med ett objekt med en blå linje i sin vänstra hand.
Barn som leker på en lekplats på en hög av däck
En man i röd snöutrustning tittar på en vidd av snö och berg.
En man som bär en hustrumisshandlare, sitter runt frukt på en låg budget marknad.
En pojke i röd hatt och svart skjorta skateboard nära en röd och vit randig trottoarkant.
Ett litet barn klättrar uppför en stenvägg i all sin skyddsutrustning.
Asiatisk kvinna i vit skjorta som står borta från folkmassan bakom henne.
En kvinna på en tunnelbana somnar.
En kvinnlig idrottsman knyter snören på en av sina klapperskor på planen.
En man i gula och gröna shorts hoppar i ett vardagsrum.
Ung flicka rör en gryta med en sked i köket medan hon bär en stor svart filt.
Flera resenärer antingen står eller sitter på vad som verkar vara en tunnelbanebil.
En pojke upplever och ställer ut på museet.
En manlig gymnast hoppar över en hög med träplattformar.
En hund travar över marken med en stor käpp i munnen.
Mannen bär skyddande ögonutrustning utför ett vetenskapligt experiment medan kvinnan klockor.
En lång man som rör om i en kruka med mat på en spis.
En kvinna blir intervjuad vid sitt matbord.
En kvinna med långt brunetthår och en beige hoodie står nära skåp.
En man med handskar jobbar i ett labb.
En pojke som ligger på gräset med en fotboll vid fötterna.
En kvinna ändrar sin strumpa i en stökig park.
Pojke och hans familj firar hans födelsedag med en ljust tänd tårta.
En man som kör ett grönt minitåg.
En man i vit t-shirt ler som om han såg på något.
En man häller drinkar vid ett bord.
Två svarta hundar travar genom ett tomt offentligt område.
En tjej i grön skjorta hoppar upp i luften.
Omkring 12 barn och några vuxna blir stänkta av en off-camera källa.
En gammal man i traditionell kostym verkar vara på ett glatt humör.
En hona med blont hår skär en vattenmelon på en marmorbänk.
Folk står på en plattform för att gå ombord på ett tåg.
En liten pojke med en blå keps sitter på en brygga med utsikt över vattnet.
Grupper av människor observerar fisk i en stor tank.
Fyra personer går över tjock snö under en solnedgång.
En servitör som lägger fram en order till kökspersonalen.
En kvinna i tölpskjorta och en beige kofta tittar bort från brädspelet hon sitter framför.
Folk väntar på sin favoritdryck.
En militär eller polis vaktar när folk passerar på ett torg.
En kvinna i röd klänning täcker en annan kvinnas ögon.
En kvinna som läser en tidning och en man i grön jacka som åker tåg.
En man som står och hejar på en stadion med andra som sitter.
En man utan skjorta går på massor av stenar.
En pojke i en röd tröja som springer på stranden
Ett par går på en sammankomst med en ballong i luften bakom sig.
En man i svart hatt går nerför gatan.
En man står på en gata och håller ett tecken.
Mannen på stranden letar efter saker med metalldetektor.
En ung pojke som bär en blå t-shirt håller upp en udda utseende objekt för inspektion medan stående bland träd.
Två små barn står i hallen.
Vattenskidåren gör en volt bakom en båt.
En liten pojke sitter på en bänk bredvid en stor geléböna maskot.
Två personer vaknar i vattnet och dras av en båt.
En man strör kryddor på sin grill framför lövverk.
Pojke med mörk hud, stående på huvudet med ben utspridda, i slutet av en flytande träbåt.
Två män spelar musik på en bänk.
Två kvinnor i färgglada kostymer tittar på en liten flicka i brun väst.
Några barn tittar på fisk i en pool.
En grävsko ligger ovanpå en hög med spillror från en riven byggnad.
Tre pojkar leker med paddlar på stranden.
En kvinna i en ljusblå jacka cyklar.
Någon tar en promenad på sin cykel.
Två personer med hjälmar cyklar framför en byggnad.
Två cyklister som rider bredvid några järnvägsspår.
Ett par njuter av en vacker dagcykling på en cykelled med bicykling skyddshjälmar och handskar.
Kvinnor i cykelhjälmar tar paus från långfärd.
En man med svart hjälm, blå jacka och khakiskjortor cyklar på gatan bredvid en röd bil.
Grabben ska åka cykel med föräldern.
Två små pojkar ser tillbaka när de går över ett gräsbevuxen område.
Barn på en liten motorcykel nära en liten damm.
Två blonda flickor i hjälm sitter på en röd ATV.
En pojke i vitt spelar baseball.
En ung pojke med tungan utstucken klättrar upp på en träplattform.
En kvinna som står vid disken vid ett takeoutfönster.
En hund med blå sele står i snö och byxor.
En kvinna står bredvid en japansk version av Disneys Snövit.
En kvinna beställer en maträtt hos en gatuköksförsäljare.
Hundar som drar en släde i ett slädlopp.
En ensam musiker i svart står på scen, spelar akustisk gitarr och sjunger in i en mikrofon.
En ung pojke i baddräkt sitter i vatten.
En kvinna i jeans går längs en stig med grönt räcke.
En kvinna i svart skjorta kramar en man.
En kvinna som hukar sig i gräset ler mot en liten pojke, när han ler och höjer händerna i luften.
Hunden har röda remmar i ryggen.
En svart hund och en vit hund står på snö.
En hund som hoppar i vattnet vid en näbb.
En brun, fluffig hund som hoppar in i en pool efter en röd leksak.
En vit hund som hoppar för att fånga en röd boll.
En pojke hoppar från ett bord till ett annat i en park.
Två och fyra fotade grannar kommer förbi för att besöka.
Ett tungt par interagerar utanför en randig cabana på en strand som ligger nära en brygga.
En ung flicka försöker ta hand om trädgårdsskötseln.
En kvinna som håller i en gul väska sitter på en stol i en affär.
En kvinna som sträcker sig ut mot ljuset.
Tre unga kvinnor uppträder en dans i en fullsatt sal.
Det finns tre simmare från samma lag som gör sig redo att tävla.
Två personer simmar i vatten bredvid en röd boj.
Två pojkar står bredvid en hög med sopor på marken.
En liten pojke håller i en grön och gul svamp medan han står framför en spis.
En kvinna som hukar sig för att möta ett litet barn medan hon håller en hund.
En man som står i ett hål framför en kvinna i en trädgård.
En arbetare i en blå hatt håller på att laga väggen.
En kvinna i traditionell islamsk dräkt går genom ett torg med en skäggig man.
En familj poserar för ett foto vid middagen.
En kvinna talar animerat med sin kamrat bredvid en vattensamling.
En man med hatt som jonglerar inför en fängslad publik.
En man på en telefon och en kvinna som sitter nära en målning.
En kvinna som håller en hund i koppel.
En person dukar vid ett bord i ett café.
En kvinna dricker av ett grönt sugrör.
En gentleman i lila halsduk och hatt tittar på pengar medan han håller i ett dragspel.
En dam i röd och svart randig skjorta sitter på en bärande vägg.
En skara människor står tillsammans på en trottoar, medan en man tar en bild.
Kvinnan i glasögon håller i en röd och vit väska.
Fyra pojkar springer nerför en stenlagd trottoar.
En kvinna tittar ut genom fönstret när en man tittar in.
En vandrare med en amerikansk flagga på ryggsäcken går genom skogen.
En man i röd skjorta sitter vid ett bord med ett glas vatten.
En man som tillagar något i en gammal brinnande ugn med ett förkläde på.
De här människorna lagar massor av mat.
En liten flicka i en tröja svängs runt av en osynlig hand.
En man i overall och hatt tenderar till en stor spole av rep.
En pojke i badbyxor gör en backflip i havet medan bergen visar sig genom dimman bakom honom.
En skadad, blodig person som sitter med vänner på ett sjukhus väntrum.
Sex skjortlösa män står utanför lutande på eller står nära ett staket.
En målare visar upp sin talang inför en grupp människor
En pojke håller i näsan och hoppar från en dykbräda baklänges in i en sjö.
En ung pojke kör en billeksak uppför en kulle.
En asiatisk kvinna i en röd tröja som håller sitt barn.
En asiatisk man ger kameran ett ont öga.
Ett litet barn som bär en sinne sträcker sig för att se ett videospel i en arkad.
En ung pojke som ligger i vattnet.
Tre pojkar i storlek för att bli blöta bredvid en vägg
En kvinna med flätor knäböjer och justerar snöret på en maskin
Två personer med gula ryggsäckar vandrar uppför en kulle.
I ett träd fyllt park en man sträcker.
Olika passagerare på en buss tittar ut genom fönstret eller in i avståndet.
Två vakter håller fast en annan man vid axlarna och armarna.
Två vandrare går nerför en torr sluttning bredvid en grön barrträd.
Pojken har blont hår och ett smutsigt ansikte.
En kvinna ser stenig ut i spegeln när hon applicerar eyeliner.
Några killar som spelar fotboll på ett plan.
En man i Hawaiisk skjorta spelar en orange elgitarr på en scen.
Människor på ett fullsatt tåg eller buss i Asien.
Det finns en man på en böljande häst som håller hårt i sig medan publiken tittar på en rodeo.
En vuxen man i jeans och svart skjorta som håller i en dryck.
En man har sina armar runt två kvinnor som poserar för en bild med honom.
En mobil matstation för att betjäna kunder på stadens gator.
En kvinna med en röd jacka och hennes följeslagare äter snacks.
En mycket ung pojke glider nerför en rutschkana i en swimmingpool och bär blå floaties.
Flicka med grön tank övredel står mitt i ett tåg spår med flerfärg tåg bilar till höger.
Tjejen står ut på tågspåren.
En fiskare förbereder sina nät inför nästa drag.
En kvinna sitter på en pall med dragspel.
Två grå hundar springer genom ett fält av rosa ljung.
En ung pojke med simglasögon, hoppar in i en simbassäng.
Folk arbetar på fabriksgolvet medan gula högar av papper går förbi.
En ung man, barfota längs stranden, beskärer ett träd.
Två barn på Wakeboards försöker ge varandra en high-five.
Ett utomhuscafé med människor som sitter medan en man i vit skjorta går mot dem.
Det finns många människor med svart hår på väg genom vissa dörrar och några kommer ut.
Flera personer går uppför en trappa.
En man klädd i en bourgogneskjorta och svarta byxor som manövrerar en marionett som håller i ett musikinstrument.
De två racers körde den vita cykeln nerför vägen.
Två pojkar, en i rött och en i vit uniform, slåss om kontroll över bollen under en fotbollsmatch.
En man i gul väst som sopar en trottoar.
En asiatisk familj lagar kött på spett på en nattmarknad.
En svart hund simmar i vattnet.
Två män, en stående och en på en cykel pratar utanför en byggnad.
Gruppen tittar på en tecknad film på en liten elektrisk enhet.
En man med en axelväska som går i öknen på sanden med fotavtryck bakom sig och horisonten med många stormiga moln.
En leende pojke springer genom gräset.
En brun häst står bakom en flicka och sniffar hennes hår.
Unga kockar ordnar mat i ett kök.
En pojke i blå skjorta som stänker i vatten under en docka
En pojke som plaskar genom havet.
Arbetare serverar kunder som står uppradade framför ett Martins berömda louisiana korvförsäljare tält
Två tjejer utför tricks på en studsmatta.
En tjej i röd bikini hoppar in i en pool.
En man drar en vagn täckt av stolar.
En hund med en röd krage och tungan som hänger ut rinner genom högt gräs.
En ung pojke som täcker ansiktet när han sitter på en studsmatta.
En leende kvinna i lila skjorta och vitt förkläde som torkar händerna på en servett.
Person som hänger upp och ner från stolpar
En man som bär en grå t-shirt och blå jeans står redo att träffa en golfboll på en driving range.
Två valpar springer över platta stenar i trädgården.
Hundar springer på en kall men solig morgon
En äldre svart kvinna kör sin elektriska rullstol.
En grön tonad hand hålls upp framför ett bord av människor.
Två män jobbar på tågspår.
En liten flicka i en utarbetad grön och orange klänning jagar en rosa och vit ballong figur.
Dessa två kvinnor har kul när de tar bilder.
En man i röd skjorta hoppar från en stor klippformation.
Flera människor rider på en berg-och dalbana medan de reagerar på att gå igenom en slinga på olika sätt.
En ung pojke undersöker ett fält av pumpor, med några redan i sin skottkärra.
Killen som spelar banjo i parken som en anka gillar musiken.
Flickan i lila topp och shorts, bär en hatt, skrattar.
Kvinnan i bikini övredelen går på stranden
En man i mörk jacka står bredvid en man klädd i brunt och sträcker sig ner i en väska.
En man på scenen framför en konsert för folk.
En glassbil stannar framför två små hyreshus.
En pojke med svarta badbyxor står i en fontän.
En ung asiatisk pojke hoppar av glädje ner i en vattenpöl, hans tunga stack ut av glädje.
Några ungar leker nära gatan.
Den här pojken leker på en lekplats med däck på.
En SCUBA dykare som simmar djupt under vattnet med en sköldpadda.
En grupp människor bär saker på en smal väg.
En brun hund sitter i ett långt gräs.
En afroamerikansk bebis kryper på golvet nära ett bord.
En man som går nerför gatan med en liten pojke.
En man bär en soptunna förbi en staty av en ängel.
En ung kvinna på en utomhusmarknad som köper bröd.
En blond tjej i vit klänning som håller en fågel i ett träd.
Två personer åker skridskor i en rink.
En liten pojke och en liten flicka ligger på en svart bänk omgiven av vuxna.
En pojke och en flicka som leker på stranden.
En äldre man bär overall och håller i en pensel.
En gammal man sover på en parkbänk.
En man med en blå keps på sover mot en sten.
En gentleman i traditionell dräkt som väver en filt på ett fält.
En man i gul skjorta dammsuger ett golv medan han tittar på kameran.
Ung afrikansk man arbetar på ett fält.
En brun hund går längs en gräsig stig med sin långa rosa tunga hängande ut.
En asiatisk man i kostym på tunnelbanan som sover.
En kvinna i vit skjorta som blandar något på köksdisken.
Människor inne i en byggnad med huvudet nedåt med utsikt utanför cyklar.
En cykelcyklist som bär röd skjorta och svarta shorts tas hand om av stadsarbetare.
En man i smutsiga jeans ovanpå en ställning.
Två kockar pratar tillsammans bakom en kaklad restaurangkalender i en tjusig restaurang.
En kvinna i ett vitt förkläde tillagar olika köttsorter på en stor grill.
En man som sitter framför en stor Calvin Klein stålreklam med ett långt instrument.
En man och en kvinna, som båda bär shorts, går nerför en trottoar.
Ett par dansare uppträder på en röd tegelgata.
En ung pojke i vit skjorta håller i ett omslag.
En man i vit t-shirt som städar upp skräp.
Äldre man i orange overall som håller en vattenslang.
2 pojkar i förgrunden i en karate tävling och tränare i bakgrunden tittar på med en annan tränare sitter vid bordet.
Individer med ballonger deltar i en promenad.
Folk som väntar på att gå över gatan framför ett apotek med upplyst skylt.
En kvinna med glas dricker kaffe på ett café.
En man i en bowlinghall som gör sig redo att kasta bowlingbollen nerför banan.
En flicka tar bort sin ögonmakeup med en öronservett.
En stor svart och vit hund springer genom ett gräsfält.
En man som studerar för sina prov utanför en bokhandel
En ung man i röd skjorta som lagar mat i en stekpanna.
En man kysser en annan man på notan och båda är i vita skjortor med svarta västar.
En grupp människor klädde sig på samma sätt när de gick nerför gatan, i en parad.
Folk står på en färgglad balkong.
Två män som slår på trummor och en man som blåser i ett horn utanför.
En bonde går sin gris nerför grusvägen.
Två tjejer i gröna stövlar och en kvinna är tillsammans.
En marknadsplats med rullande vagnar som säljer frukt.
En kvinna med blont hår och solglasögon som sitter vid ett bord och ler.
Tre arbetarklass afroamerikanska män är utanför.
En liten flicka svingar i en baby sving på lekplatsen.
En flicka som står i havet
Två barn är på stranden och leker i den våta sanden.
En ung kvinna som ler på avstånd njuter av ett bubbelbad.
Ett barn som bär svartvit badutrustning knäböjer i grunt vatten över en plastgul båt fylld med våt sand.
En man breakdansar på golvet runt en massa människor.
En man och kvinna njuter av en tur nerför forsarna en varm dag.
En flicka som gör ett delat handstånd på stranden under dagen med en nöjespark i bakgrunden.
En man i orange skjorta använder en scraper i en sifter.
Två tjejer sparring med en röd och blå fladdermus medan en annan flicka tittar.
En kvinna knuffar en ung flicka i en gunga.
Två pojkar poserar i blå skjortor och khaki shorts.
En grupp människor väntar på en plattform medan ett tåg passerar dem.
En liten flicka som leker, på trottoaren, med en pinne.
En man som trycker på en handtruck med lådor böjer sig över för att plocka upp ett päron.
En försäljare som står i fönstret i sin butik.
Flera män av indiskt ursprung samtalar, och i synnerhet en av dem verkar mycket entusiastisk över samtalet.
Ökvinna som lagar mat utomhus med ananas och frukt.
En grupp människor i kilts spelar musik medan en löpare i svart springer förbi.
En man som öppnar en grillugn medan han håller i tången.
Den lilla flickan bär en denimklänning och håller i en brun nallebjörn.
En man fångar en hyfsad fisk och tar av den från kroken
En man med en hästsvans och solbränna som sitter på en soffa och räknar med fingrarna.
En man med grön skjorta på fungerar.
Två unga attraktiva kvinnor med shorts korsar en gata i en livlig stad.
Mannen klättrar genom klipporna och snön.
Den här bilden är av en ung flicka som tränar gymnastik i ett gym.
Två beige hundar leker i snön.
En man som håller på att kliva av kanten av en ökenstensformation.
Tre kvinnor i klänningar och huvuddukar utanför.
En liten pojke och hans cykel sitter utanför Kuthhoop Hotel.
Solen bakom en grupp träd på en lång ridning.
En man i orange skjorta tar en bild.
En publik hejar på ett baseballlag.
En man och en mycket yngre pojke, båda klädda i hattar, tar en promenad genom naturen.
En liten pojke knuffar upp en pojke till.
En man med vit skjorta och slips står på en trottoar mellan cementbarriärer.
En pojke når toppen av ett djungelgym.
Två personer i svarta västar står framför barn i vita västar med en amerikansk flagga mellan sig.
En man med svärd som slåss mot en kvinna med ett spjut.
Två män mitt i en match.
En ung man i en vit skjorta som skär tomater.
En ung pojke i blå shorts klättrar klippor längs hotellet resort strand strand.
En man spelar saxofon bredvid en gul brandpost.
En man på fiskmarknaden skär svärdfisk till stekar.
En hund i luften som tar den röda bollen.
Tre kvinnor klädda i vanliga kläder lagar mat i köket.
Folk går och springer på en trottoar.
Två unga kvinnor går längs en landsväg som gränsar till träd.
En ung flicka på stranden som springer mot vattnet.
En ung pojke i blå skjorta och grön hatt spränger en orange ballong.
En svart och vit hund som hoppar in i en pool efter tennisbollar.
Den lille pojken springer åt fel håll efter att ha slagit bollen i en omgång tee-boll.
En person i en blå skjorta håller en mikrofon i sina händer.
En man i vitt och rött med solglasögon som bär och blåser ett mycket stort horn.
En rödhårig barfota flicka som hoppar över en rail.
En kvinna i shorts kastar en bowlingboll i en bowlinghall.
Han läser en tidning och hon tittar på honom med ett leende.
En brun hund på ett koppel som springer i grunt havsvatten.
Pojken hoppar i skogen.
En man och en kvinna sitter på marken och omges av båtar.
En ung pojke på stranden som springer in i havsvågorna.
En pojke i en blå båt som är fastbunden vid en större båt dumpar en hink vatten.
En man som går på en smal gata.
En ung man vilar på en flygplatsplats med en cowboyhatt över ansiktet.
Barn som fiskar vid en bro
Man sitter i skuggorna på trappan i en byggnad.
En svart och vit hund som hoppar in i en pool.
En svart hund och en vit hund ras i ett gräsfält medan åskådare tittar på.
Ett gäng fåglar utanför en byggnad.
En golfare förbereder sig för att ta ett skott på golfbanan omgiven av träd.
En brandman släcker en brand under motorhuven på en bil.
Folk samlas runt ett bord med många röda, vita och blå dekorationer runt i det rymliga tältet.
Ett litet barn med ägg i en skål.
Tre tonåringar bär ved på en gata medan en av tonåringarna ler mot kameran.
En man står framför Gateway Arch.
En ung pojke med bläck står framför en vit dörr.
En blond tjej trampar på vertikala stockar i sanden.
En ung flicka med lila skjorta, vattengräs.
Katten ser bort från personen bredvid.
Ett par väntar på en korsning i en ljust upplyst stad.
En person i gul skjorta som sträcker sig på en bro.
En magkänsla med en rutig skjorta med mustasch som säljer fisk på en marknad.
Stadsarbetare gör underhåll på en tågbana.
Ett barn framför sin egen spegelbild vänder sig mot kameran och ler.
Arbetare lastar funktionshindrad man i rullstol på ett tåg.
En kvinna som går på en gata med en ung pojke framför sig, och en löpare bakom henne.
En kvinna ser upprörd ut när hon håller en vattenflaska framför en vägg och skriver på den.
En grupp afrikanska pojkar tittar på vattenledningar.
Tre människor på gräs, en krattande löv, en klippning gräsmattan, en annan stående vid en soppåse.
En pojke med gul skjorta och svarta byxor som svetsar något.
En man utan tröja klättrar på en sten.
En tjej är på väg att kasta en softball.
En man kastar upp ett litet barn i luften.
En fluffig vit hund kommer ut ur en blå randig hindersluss.
Två barn sitter på golvet tillsammans.
Ung flicka bär campingutrustning och en uppstoppad brun hund.
En kille med grön skjorta lagar mat på en lägereld.
En flicka kikar genom löven på ett träd.
En motorcyklist kör upp på sidan av ett grönt berg medan en annan cykel förblir stationär.
Ung pojke i klättring sele skala en klättervägg.
En man vadar i vattnet och tittar på ett vattenfall.
En svart hund går genom en ström av vatten.
En man surfar nerför en sandkulle.
En man med röd-rimmade glasögon står med armarna vikta bakom en metallgaller.
En hund springer medan han håller ett föremål i munnen.
En hund med långt hår och en röd väst går i gräset.
Två poliser i uniform som chattar i en golfvagn.
Yngre man i gul skjorta och bruna shorts flyttar en torr gård eller åker med en ridning John Deere traktor flyttare.
Säkerhetsvakten ler.
En lång dag gör kvinnan trött och sömnig.
Vacker brunett kvinna, dragen i lila, blå och en scharlakansröd scarves.
En liten svart hund är i gräset.
En flicka i en grå YMCA-tröja tittar genom ett teleskop.
Ett barn försiktigt insvept i en filt som sover i en sjuksäng.
En ung dam som spelar gitarr på en scen i en park.
Tre små pojkar tar ett bad i en gummibehållare på gräset.
Flera personer sitter vid datordiskarna på ett rörigt kontor.
Flicka med halv dreadlocks och öronmuffs på gör en stor bubbla
Barn och kvinnor samlas utanför en byggnad.
En man kryper genom en lekplats plaströr mot en liten flicka med rött hår.
En flintskallig man klappar en vit panda i ett zoo.
En skjortlös man i blå hatt och solglasögon löper midjedjup genom en stor vattenförekomst.
En man i svart skjorta och hatt spelar gitarr.
En man i vit skjorta plöjer ett fält med två mulor.
Folk som leker i vattnet med en vattencykel.
En blond person rider en jetski i vatten nära en bergskedja.
Två man sitter i vitt rum och spelar gitarr.
Tre kvinnor går tillsammans längs trottoaren, en bär en kort vit kjol.
En pojke håller händerna på huvudet.
En man målar stänkta kläder talar på en mobiltelefon.
En man i fönstret på en röd lastbil.
En man i orange regnrock diskuterar något med en annan man som bär arbetskläder nära ett kloakhål.
En man i svart skjorta står framför en byggkon.
S stor man i en blå skjorta och shorts lutande mot en van framför en butik som heter "Terrible's"
En videoograf och en kvinnlig följeslagare står vid en vattenväg.
En regnbåge bildas av en tank som sprutar vatten på en gata.
Mannen med bockskjorta och svart skjorta går längs gatan.
En man i grå skjorta och en hatt som håller en jackhammer
Två byggnadsarbetare pratar när de tittar på ett marinskepp.
En person som hoppar från en sten på en smutscykel.
En tjej som spelar pool i en poolhall.
En man klättrar uppför en klippa och når ett överhäng.
En grupp människor som går över en repbro.
En ung man ensam på en vitsandsstrand har ett mellanmål under ett strandparasoll.
En man uppträder för en publik på en lång enhjuling.
En ung pojke springer nerför ett fält och bär en namnbricka.
Jord, vatten och himmel gör detta till en bra plats en timeout.
Ett ungt barn som bär blå sovkläder har en napp i munnen och sover.
En man och kvinna går längs gatan tillsammans.
En kvinna ler och läser en tidning bakom en lätt reklam.
Två personer tittar över en terrassvägg.
En kvinna med motorhuv sitter ner med händerna i knät.
Tre arbetare arbetar på ett metalltak
En kvinna med slitna jeans ligger på marken med underarmen över ansiktet.
Kvinnan går med ansiktet målade barn medan bär ett skrikande barn.
En kock med glasögon lagar franskt bröd i en jätteugn.
Två personer står utanför en vinbutik.
En man och en kvinna tar sig utanför ett kaffehus.
En silhuett av ett barn som leker på en strand.
En man med shorts, sandaler och en svart skjorta pratar på sin mobiltelefon.
Två män pratar i ett restaurangkök.
En ung flicka sitter på en klippa med utsikt över ett stort fält.
En man i grön hatt som springer.
Två hanar springer, en bär rött och vitt, den andra marinblå och svart, utanför en molnig dag.
En liten pojke i gul skjorta som går på stenar.
En skara män och kvinnor som står och står vid en vi kräver tecken.
Fem asiatiska vänner poserar tillsammans för en bild.
Fyra kvinnor och en man sitter på trottoaren med sovsäckar.
Många människor samlade ihop
Tre ungdomar smyger under en filt på en trottoar.
Två personer tar bilder.
Tre kvinnor och en man i en hatt sitter korsbent i en grupp.
Det är en asiatisk flicka som har en grön skylt som protesterar.
En man som filmar en grupp människor framför en New York-banner.
Människor på en gårdsplats sitter och står.
En man i limegrön skjorta väntar på tunnelbanan medan en kvinna filmar med sin telefon.
Unga människor i gula skjortor tillagar färgstark mat.
En kvinna i gul skjorta hjälper en liten flicka i rosa skjorta.
Ungar serveras gröna ägg och skinka.
En man i en blå skjorta som håller ett barn medan han håller i en barnvagn på en basebollstadion.
Små pojkar i vita karate uniformer utför sina kampsporter inomhus.
TVÅ människor går in i en skugga i en riktning medan en annan går mitt i den.
En man, en kvinna med barn i en barnvagn på en fullsatt gata.
Mannen siktar på att skjuta något medan hans hund tittar.
En häst går bredvid en båt under en bro.
En ung man sitter vid ett bord med en laptop och hörlurar.
En man spelar banjo på en konsert.
En dam med en väska tittar på varor på en loppmarknad.
En man åker snowboard över en byggnad på en snöig kulle.
Den bruna hunden ligger på ett blått lakan.
En man i svart skjorta som läser en tidning.
En man som bär glasögon och en blå jacka ler medan män bakom honom lagar mat på en grill.
En kille i skinnjacka som går förbi en hörnbutik.
En grupp vänner står framför konsten de har sprejat för en bild.
Han gör stunts med sin cykel.
En kvinna tittar på klädda, huvudlösa skyltdockor i en butiksutställning.
Ett barn som står mitt på en grusväg
En man i brun skjorta tar en bild av något på marken framför sig.
Folk som sitter framför andra människor.
En man som bär en brun t-shirt pratar med en kvinna som bär en blommande tanktopp på en utomhusmusikkonsert.
Två flickor på stranden tittar på folk i en båtfisk.
Två cyklar står bakom två personer som sitter på gräset nära en vattenförekomst.
Två gamla män sitter på bryggan.
En man i kostym och två män i orange väst.
Ett litet barn knuffar en barnvagn nerför gatan.
En kvinna vid examen utan mössa.
En äldste man har utsikt över en balkong som vetter mot en gata.
Den här kvinnan ler och pratar i telefon medan hon sitter på en stenvägg.
Tre hundar på ett fält tittar på något i gräset.
Tre barn, två flickor och en pojke, i kampsport ställning, står på hårt trägolv i ett stort rum.
En kvinna sitter på en blomkruka på ett fullsatt kafé.
En pojke står bredvid ett räcke vid en go kartbana.
En vit fågel står på en träplattform.
Det är en kille med styltor som spelar trombon framför en väggmålning.
Två unga pojkar, som bara har underkläder, klättrar runt ett fordon.
En ung blond tjej i rosa skjorta tittar på en stor bönemantis på armen.
En man klädd i vitt och med glasögon som har något att äta.
En man fiskar längs en strand i en stor vattensamling medan en ung pojke bär ett nät inte alltför långt bort.
Soldaten står lång när han ser det förbipasserande folket.
En ung man i kostym står ut från publiken, på vad som verkar vara en konstutställning.
En man som bereder frukt under ett träd.
En svart hund kommer ut ur havsvattnet på stranden med något i munnen.
Två små barn leker på stranden medan en man tittar.
En grupp människor sitter på en strand och tittar på Blue Angels.
Två unga damer spelar schack på en restaurang.
En person som bär en långärmad vit skjorta väver med gul tråd.
Två kvinnor joggar och tre män går på en grusstig.
Dessa är kvinnliga medlemmar av en musiksymfoni klädd i svart och bär röda flaggor utanför en utsmyckad byggnad.
En familj på fyra tittar på en flygshow.
En person som håller en liten hund i koppel böjer sig över och tittar igenom föremål.
En brun hund som bär på ett svart föremål.
En rädd liten pojke som dras upp och ur en pool av sin far.
En man som står framför flera klippor.
Två personer och en liten vit hund leker i parken.
Två män med långt hår sitter på marken.
Medlemmar i ett mässingsband tittar på sin noter.
En man spelar ett DJ-spel i en arkad.
En grupp kvinnor klädda i svart spelar musikinstrument framför en stor byggnad.
En man sitter ovanpå en skolbuss, medan en annan man, som bär en matchande skjorta, står inne.
Demonstranter som väntar på att polisen ska höra deras klagomål mot polisförtryck och brutalitet.
En man som bär cowboyhatt och ett guldkors runt halsen
En gammal man och en ungdom jobbar på att starta en ror.
Folk väntar på sitt bagage på flygplatsen.
En grupp människor utanför efter mörkret mot en vattenväg.
Fyra kvinnor deltar i synkroniserad simning i mörkret.
En brun hund jagar en blond i gräset.
En man i svart hatt och solbränd jacka som går tvärs över gatan.
En ung flicka som bär bikini i ett innerrör.
En man som bär långt hår syr en kostym.
En man med brun t-shirt håller i en tråd medan en annan man tittar på.
En man i en mantel är nära en röd byggnad.
Två män klädda i business casual dela ett skratt.
En basist i röd skjorta spelar medan man röker en cigarett.
En svartklädd man med udda huvudbonader svänger en stav.
En mager flicka i stora stövlar står vid vägkanten.
Två kvinnor står på en båt och tittar på vattnet.
Folk tittar på bilder på en display.
Den lilla flickan sitter i en sele, fastspänd i en tjuder, medan andra tittar.
En man som bär en mångfärgad skjorta håller i en megafon.
En ung man med mörkt hår och skäggkokande biffar ute på en liten grill.
En uniformerad kvinna som håller en kamera stående framför en skara åskådare.
Den lilla pojken i röda trunks försöker fånga en fotboll som kommer mot honom.
Fyra ungar rullar och glider ner för en sanddyn.
Den lilla lurviga vita hunden går i det gröna gräset.
En liten flicka high-five är en gul robot.
En person klädd i en blå skjorta och jeans ser förbi träden till horisonten.
Gråa och svarta hundar springer iväg längs skogsstigen
En kvinna och en ung man dukar vid ett bord i en mexikansk restaurang.
En bergsklättrare stiger upp.
En dam i svart klänning pratar med en grupp människor.
Två män sitter och jobbar på sina datorer.
En man som häller en skottkärra cement på en trottoar.
En hund springer längs den korta på en strand.
En ung gentlemän med en blå slips som pratar in i en mikrofon.
Flera yngre människor går nerför en gata i tunga kläder.
Kvinnor av olika etnicitet står i ett rum, håller röda och gula pilar.
Två hundar skakar av sig vattendroppar på en strand.
Den manliga bergsbestigaren tar en titt över axeln på utsikten över sjön och staden.
En man som klättrar tar en paus för att beräkna sin rutt.
En brud och brudgummen matar varandra med bröllopstårta.
Fem arbetare som sitter framför lastbilar och äter lunch
Ett ungt gossebarn med lockigt brunt hår, som gömmer sig bakom en kartong på en grönsaksmarknad.
En kvinna ligger i gräset och äter något utanför pizzatornet.
En man och en kvinna spelar på ett kasino och roar sig.
Skäggig man som spelar akustisk gitarr
Ett barn lyckas dra sig till fötterna med hjälp av en soffa.
En man arbetar på en träbit på en spinnare.
En man med säkerhetsutrustning driver en maskin med tält på bakgrunden.
En kvinna, klädd i gul blus och svarta trosor, spelar beachvolleyboll.
En flicka ler när hon springer över den vita sandstranden i baddräkten.
En man i svart skjorta hoppar med en kaffekopp full av en dryck.
En man som leder en KitchenAid-klass klädd i en svart kockjacka.
En man skålar med sin drink.
Mannen i en mörkblå skjorta kramar en flaska fylld med ett guldfärgat ämne.
Folk i en affär utanför under ett tält.
En grupp damer med datorer sitter bakom ett bord medan folk på andra sidan köper något.
En man i en vit kockjacka med tomater.
En kock pratar med en annan person i ett KitchenAid showroom.
Många människor samlas under ett tält och får mat.
Ett barn står på sidan av en soffa och slår över en lampa.
Mor och far ser på när deras barn klappar ett djur.
En man arbetar på en mycket stor, invecklad sandskulptur på en strand.
Tre personer sover i en masstransitbil.
En man i jacka, hatt och huva, vänd mot kameran håller händerna upp och samman.
En man och en kvinna med shorts står i en gränd.
En pojke gungar ett basebollträ, och en fångare står bakom honom.
Två små ligor är bredvid en bas på fältet.
En ung man med blont hår arbetar med flerfärgade trådar medan han sitter på en stolpe.
En kvinna i svart jacka lutar sig mot en lyktstolpe.
En mörkhårig kvinna i svart skjorta tittar på en silvermaskin.
Två kvinnor och ett barn i en barnvagn framför en affär.
En man i randig skjorta spelar trummor.
En person som ser ut och står på en sten.
Ett barn hoppar på en sanddyn.
Två tjejer som sitter vid vattnet.
En ung pojke står i ett klassrum och försöker göra ett pysselprojekt, men har svårigheter, medan hans klasskamrater tittar på honom.
Två dansare på scen i en klubb.
En gentleman skrattar i sin bil när han kör på landsbygden.
Tre pojkar krossar tegelstenar i små bitar.
En man i en färgglad skjorta och en dam i en vit blus signerar böcker för människor.
Tre kockar lagar mat i köket.
Fem kockar står bakom ett bord fullt av muffins.
Män och kvinnor och Michigan Vin- och matprovning
En pojke leker med utsträckta armar på trottoaren bredvid en kullerstensgata.
En man i röda badbyxor som spelar volleyboll.
En äldre dam i svart skjorta är att lägga ingredienser till en KitchenAid blandning skål som en publik ser på.
Folk sitter på barer med en massa vinglas.
Ett sportlag som består av 14 kvinnor med vit t-shirt och rosa taggar.
En kock som lagar hamburgare utanför, på en grill för gäster som går förbi.
En ung pojke i Tigerskjorta står ovanpå någon som ligger i en säng.
Två män jobbar på taket av en byggnad.
Folk är på en åktur som sänker en från en hög höjd.
Man i svart på mikrofon, i band.
En man och en kvinna går i en äppelträdgård medan de svingar en liten pojke mellan sig.
Den unge mannen håller ett glas och kollar sin mobil.
Två små pojkar sitter i en metallformad låda medan de bär cykelhjälmar.
En grupp människor som verkar ha roligt.
En kvinna i röd träningsoverall som klämmer citroner i en press.
Flicka och pojke serverar mat på tallrik
Två barn med brunt hår i bakluckan på en bil.
Ett litet barn håller huvudet av sin äldre bror
En man som bär vit skjorta och handskar håller i en rutig låda.
Street scen i Asien med fotgängare och parkerade cyklar.
En våt hund hoppar över ett hinder.
En kvinna tar tag i en killes fot och lägger den bakom hans huvud.
En kvinna, i nunnekläder, blir friterad av en kvinnlig säkerhetsvakt, medan en annan kvinna tittar på.
Mannen i mörk kostym håller på med en pratradioshow.
En fiskare rullar sitt spö medan en annan slappnar av i en båt på vatten.
Folk samlas utanför för en protest, och en kvinna längst fram ler mot kameran.
Personen bär en svart och röd dräkt och övar strid.
Ett barn i en ninja outfit gör en hoppspark.
En ung flicka flyttar några resväskor som är nära ett öppet fönster.
Folk sitter och ligger på trappan.
En man i vit skjorta som spelar en svartvit gitarr.
En man bredvid en clown med andra människor i bakgrunden.
En äldre dam blåser ut en 9 och en 0 nummer ljus på en födelsedagstårta.
Handyman arbetar på ytterväggen i stadshuset.
En man i gul jacka tar en bild medan han lutar sig mot en bil medan en annan man arbetar på bilen på motsatt sida.
Två personer äter en måltid tillsammans.
En man på ett fält bär ryggsäck och det finns får och berg bakom honom.
Tre brandmän samtalar bredvid en brandbil.
En stadsmarknad på en gata ligger i förgrunden, med stadsbyggnader låg i bakgrunden.
Vissa människor är på en uteplats och det finns en brand.
En man sitter på ett fält nära en ryggsäck.
Byggarbetare som arbetar på en stor byggnad.
Två leende små blonda tjejer i rosa byxor svingar från en metall bar.
Lilla pojke som går med käpp på spår
Två stora schäferhundar leker i vattnet.
Hunden hoppar i luften för att fånga en boll.
En liten flicka klädd i gult håller i två röda handtag.
En blond tjej som sitter med ett barn.
En unge i blå jeans och svarta strumpor sover under en rosa filt med en virveldesign.
En man i vit skjorta borstar en get.
En flicka med slutna ögon rör vid en pojkes kinder.
En man i vit skjorta balanserar på vattenfyllda tankar som innehåller krabbor och fisk.
En grupp människor sitter och tittar på en händelse bakom en Tim Hortons skylt.
En man står och läser något genom ett räcke med utsikt över en stad.
En ung pojke med blomma i ansiktet blandar deg i randig skjorta, overall och förkläde.
En ung pojke håller i ett blått handtag på en pier.
En man talar in i en mikrofon, medan en annan man funderar över situationen.
En man sover ute på kartong bredvid en vattenflaska.
En liten flicka klädd i en vit klänning förbereder sig för att lägga blombladen ner för ett bröllop.
En åkare rider sin bräda på en ramp.
En man i shorts står på en stol och gör en hydda.
Två vandrare som bär mörka kläder vilar på en snötäckt topp.
En man med utsträckta örsnibbar med svart hatt står framför en uppvisning av mat till salu.
En man som fiskar vid en brygga vid solnedgången.
En man klättrar på några metallstavar som är fästa vid varandra.
En liten unge som sitter i en traktorklo och leker i smuts.
En vit hund med en pinne i munnen som står bredvid en svart hund.
Paret kysser varandra, medan de står ansikte mot ansikte.
En man med röd hatt och en penna bakom örat ser ut som om han är på väg att säga något.
En ung dam som bär gul matar ett litet barn vid bordet.
En man med gul skyddsväst och hård hatt kör en traktor.
Människan står utanför mot väggen med tennisracket i mörker.
Två kvinnliga beach volleybollspelare, vända mot varandra, förbereda sig för att slå bollen.
En man håller en fisk i båda händerna.
En man som bär glasögon tittar på ett runt spegel objekt hängande uppifrån.
Fem åskådare tittar på två bilar som tävlar på en kapplöpningsbana.
Flera personer sitter på filtar i en park med blommande rosa körsbärsblommor.
En man på scenen som spelar gitarr.
En vandrare går en trädlös stig uppför en kulle.
Folk står nära en matförsäljare i en park.
En man med baseballhandske är på ett fält som lutar sig åt hans sida.
En sous-chef hackar en gurka för en sallad.
Det ser ut som om de listar ut namn, för vad som finns i flaskorna.
Det finns många olika färgade bollar.
Hunden vadar genom grunt vatten och håller något i munnen.
En man i gula byxor uppträder för en publik.
En ung man i gula byxor dansar medan en skara tittar på honom.
Person med ryggsäck i fält
En liten grupp människor sitter på stranden av en stor vattensamling i gräset.
En man som stirrar in i kameran när han skär citroner.
En grupp ungdomar står och sitter runt ett bord och äter och dricker med varandra.
En asiatisk kvinna som äter med en sked.
En man i orange skjorta hoppar medan han spelar en stor trumma.
En kvinna med glas som dricker ur ett glas
På en gatufestival lagar en pojke och en man något slags "Texas Smoked" kött medan fotgängare passerar förbi.
En äldre och yngre man skakar hand på en basketplan.
En vit man med hår och skägg med ett barn på axlarna.
En man faller från taket på en säng.
Ett litet barn håller en mopp bredvid en tvättmaskin och torktumlare.
En vandrare som kopplar av på en lersluttning.
Tre killar grillar på en grill på en veranda med ett vitt staket.
Blond kvinna som ligger på en soffa och putsar läpparna.
Man på motorcykel ridning i torra fält med hjälm och ryggsäck
En person är smutscykling över klippor och vatten.
Två små barn leker med stora hjul i ett urbant område.
En kvinna i vattnet slår en säck i en sten.
En taxi med en mamma Mia-annons ovanpå.
Den vita hunden med svarta fläckar fångar en röd frisbee.
En person hänger på en klippa när de försöker klättra.
En person som klättrar på en stor mosstäckt klippa
En person står på toppen av en klippa med utsikt över land.
En man klättrar upp för en klippa.
En man som klättrar i skogen omgiven av ljus.
Ett lyckligt par som njuter av sitt utomhusbröllop.
En ung pojke slår en boll av en tee.
En man i gul skjorta som tittar ner på marken.
En man hoppar i luften framför en kustscen med vatten och berg i bakgrunden.
Två hundar i vattnet slåss om en pinne.
En trefärgad hund hoppar och fångar en rosa frisbeen som en man i shorts har kastat.
En grupp killar samlades och drack på en bar.
Byggarbetare mitt i arbetet med ett hus.
En man sätter upp en stege i ett rum.
En grupp människor tittar på en fontän i en stads skyline med palmer.
Små barn, som alla sträcker sig runt ett osynligt föremål.
En liten flicka som försöker vara som spindelman.
Ung flicka glider nerför en uppblåst rutschkana
En man och hans fru går hand i hand nerför gatan.
Två unga pojkar springer vid vattenbrynet.
En hund märker en tupplur på en matta nära sin favoritleksak, en plyschcentiped.
Chevrolet bil som visas på en sammankomst
En grå hund klättrar upp för en låg trädgren i en park.
Två flickor leker på en inhägnad ute på fältet.
En ung brun valp drar en lummig gren i tänderna på en bakgård.
En man som njuter av sitt hantverk av träbearbetning.
En kvinna visar upp en nybakad paj genom att hålla den över huvudet.
En kvinna med höga klackar och hatt.
En kvinna svänger på ett rep med utsikt över ett rött bondgårdshus och gated betesmarker och höga träd.
En ung pojke med glasögon paddlar kajak i lugna vatten nära ett stort träd.
En Jack Russell Terrier mäts för distanshoppning när han försöker fånga en frisbee.
En kvinna i en blå skjorta som gör keramik.
Två unga pojkar som springer på ett gräsfält
Två hundar leker på ett gräsfält.
En flicka tar en bild med handen över kameralinsen.
En man sprutar en design i sand
Två personer i föråldrade kläder poserar framför en snabbmatsdisk.
Två skrattande kvinnor sitter vid ett bord med drinkar.
Två arbetare är på en körsbärsplockare, den ena lutar sig ut med en säkerhetssele och den andra ler mot kameran.
Man i hatt och rock läsa tidningen nära soptunnor och graffiti.
Folk passerar varandra på en livlig gata medan de pratar på sina mobiler.
En flicka med grissvans ler.
En pojke sitter i en leksaksbil medan han dricker ur sin pipiga kopp.
En tekniker böjd över att fixa en maskin.
En man i orange skjorta står bredvid en maskin
En man i formella kläder spelar gitarr och sjunger.
En man som lagar eld i fem krukor på samma gång!
Två pojkar gör löjliga poser bredvid ett tecken.
Nygift man och kvinna hoppar av glädje på kinesiska muren.
Det finns en asiatisk kvinna som står nära korgar fulla av apelsinfrukt.
Två kvinnor ligger upp och ner på en vit säng.
En man kör en blå gaffeltruck genom en folksamling.
En man i vit t-shirt utför tricks med en jojo.
En ung man tittar inuti munnen på en ödla som figur.
Två män sitter bredvid varandra på vattnet i en båt.
Två baseballspelare står vid kannan och viskar till varandra.
En stor svart hund jagar en stor brun hund med ett grönt föremål i munnen medan en annan stor brun hund taggar bakom.
Fyra tjejer poserar framför en publik.
En gammal man i grön skjorta sitter på trottoarkanten och håller i en kamera.
Damen i tryckklänningen strippar mat till middag.
En liten pojke gör ett hjul på stranden.
En man med getdjur rider en rulltrappa.
Ett barn i en blå mössa är nära ett omålat trästängsel.
En vit man som tar en promenad.
En egret står på en klippa vid kanten av en flod.
Man paddlar i blå kajak i vattnet.
Den skoputsande mannen, som försörjer sig på skor, skiner på en mans svarta läderskor i fina klänningsbyxor.
En man gräver ben och verktyg från en arkeologisk plats.
En grupp män står runt och dricker vatten med sina cyklar.
En afrikansk pojke kör sitt team av oxar på en grusväg.
En man spelar gitarr i en park medan folk sitter på bänkar.
Den feta, gamle mannen somnar i stolen.
En man i vit t-shirt håller paraply och glass vagn.
En man i jeans och en grå skjorta som står bakom en sprejmålad tegelvägg.
En flicka i randig skjorta håller en bulle i munnen.
Fem personer spelar stränginstrument offentligt.
En person i brun skjorta knuffar ett barn i en barnvagn vid havet.
Två personer som försörjer sig på kläder och lagar mat på ett berg.
Tre män i fiskemössor står på klippor.
Den barfota kvinnan i solglasögon sitter i trädet.
En grupp människor går på en stig nära sjön.
En man i grått håller hundens koppel medan hans son sitter på axlarna.
En man sitter i ett rum bestående av träpaneler.
Fyra tonåringar i skoluniform går längs en tropisk väg.
En ung flicka med målat ansikte står bredvid några andra barn.
Två kvinnor rider sina trehjulingar.
Den svarta hunden och den vita hunden verkar vara redo att slåss.
En gitarrist spelar medan folk leker med hula-hoops i bakgrunden.
En ung pojke bär en röd halsduk runt huvudet med ordet fri skrivet i rött på ena kinden.
En dam i blå klänning som sjunger.
En sångare och hennes band uppträder på scen i en klubb.
En man som spelar gitarr med sitt band
En man en kvinna och ett barn sitter på en soffa leende
En ung flicka hängd med rep bredvid ett nät.
Tjejen i blå jeans och vit skjorta balanserar på ett ben.
En pojke på en lekplats gunga slår en medatativ pose.
En man som bär en grön nummer tjugofem jersey sparkar en vit fotboll på ett fält.
En man rör vid sidan av ansiktet.
En liten pojke står bredvid ett fönster och gråter.
En man städar sin båt på uppfarten.
En man i grön skjorta och brunmössa lutar sig mot ett räcke i någons kök.
En kvinna som röker en cigarett lutar sig över att prata med någon.
En svart man sitter uppmärksamt vid sin symaskin omgiven av färgstarka tyger som hänger på utsidan av en succobyggnad.
En man som sitter utomhus stryker tyg medan tre personer observerar
Två unga flickor sitter i vardagsrummet och spelar TV-spel och dricker läsk på burk.
En liten pojke försöker laga sin cykel.
Den svarta hunden kommer fram ur vattnet efter att ha samlat ett föremål i tänderna.
En man med en röd hjälmkajak.
En man i kajak som simmar i grova vatten.
En person i en skyddsväst som knuffar en lastbil.
Tre män i orange västar drar en jeep ur en ravin medan en annan man sitter inne.
Två män med vita cowboyhattar.
En brun hund springer genom gräset och håller något i munnen.
Få damer går barfota på stranden.
En man som bär flytväst använder en karta på en liten båt.
Två unga flickor bär rosa spel på en lekplats
En man i vit skjorta spelar gitarr för en kvinna i vit skjorta.
En baseballsmet som lyfter armen.
Kvinnor som bär föremål på huvudet går längs en grusväg med grönska på varje sida.
Två tjejer på ett djungelgym.
Han har säkerhetsutrustning på sig medan han tränar den svarta hunden.
En man som bär färgglada kläder och vita solglasögon spelar en stor trumma med händerna.
En ung pojke i en pool som leker med en grön vattenpistol
Brun hund ligger på grus med gräs och träd i bakgrunden.
En portal man i orange overall står bredvid en grå kvinna på motorvägen med en motorcykel på sidan mitt på motorvägen.
En man som kör traktor drar med sig två små barn för en åktur.
Två personer går ut i ett naturområde.
En man och hans hund i bergen.
Två pojkar går in i en skåpbil och en yngre pojke sitter i en bilstol.
En grupp barn som leker med däck.
En kvinna som sitter på tunnelbanan håller i en vit låda medan hon blundar.
Två hundar leker med varandra
En svart hund som springer ner i vattnet.
En liten hund och en stor hund med ett rep i munnen.
En man i kostym går förbi en byggnad medan motorhuven på en bil speglar en förvrängd syn på den byggnaden.
Person med två skidstavar som åker nerför en snöig kulle.
Sju personer rider en grön flotte i en vitvattensälv.
Många går genom en park med många träd.
Kvinna i vit topp och gröna byxor som hanterar gröna grönsaker.
En man går tvärs över gatan.
En stor kvinna med kort hår som sover i en stol offentligt.
Människor går runt i en nattlig miljö.
En man skär upp mat för att lägga i skålar med mat på en matgård.
Fyra skidåkare som klättrar på snötäckta berg.
En ung flicka med blont hår och glasögon sitter vid ett bord i en restaurang.
En person forsränning i turbulent vatten.
En ung man i shorts tittar in i en bäck bredvid en klippvägg.
En pojke på en grön plastsving.
En man i blå skjorta är på väg att korsa gatan medan en polisbil kör förbi.
Den lille pojken leker med däck.
En kvinna som äter lite mat medan hon sitter på en liten pall bredvid en propangrill.
Kvinnan i blå shorts går barfota på stranden
Två män i teal scrub står framför ett café med en öppen skylt.
En person i en kilt går längs en överfart.
En pojke och en liten pojke står vid en vattenfontän.
En grupp människor går till stranden.
En surfbräda som dyker upp ur havet med sin bräda, när vågorna rasar i land bakom honom.
Fem ungdomar lagar mat i ett kök medan de tittar på TV.
En ensam bergsklättrare i en sele klättrar på en stor bergvägg.
Närbild av mannens ben på en cykelpeddal.
Fem män tvättar fönster i alpina byggnader på fem stegar.
Folk klättrar upp i en egendomlig barrerad byggnad.
Brun och vit hund som springer genom höstlöv på marken.
En pojke skateboards och gör ett hopp över en annan skateboard.
Ett lerigt barn hoppar ner i mer lera på marken.
En kvinna i grön jacka trycker på knappen för att korsa gatan.
Ett äldre par går förbi en juvelaffär en solig dag.
En smal bäck löper mellan lövtäckta kullar.
En man i dykardräkt har en låda.
En tjej på stranden som precis kom ut ur havet.
En ung man som håller en ölflaska och en cigarett stänker vätska på kol i en grill.
En flicka som ligger vid gräset
Scuba dykare under vattnet håller små kräftdjur i sina händer.
En liten flicka som springer nerför en upplyst korridor.
Unga asiatiska flickor vilar längs flodkanten.
Tre personer poserar framför en stor vit byggnad.
Unga studenter spelar musikinstrument i en orkester.
Två män är under jorden och verkar vara gruvarbetare.
En mörkhyad man i en halmhatt som spelar gitarr och en man i solglasögon som lyssnar och ler.
Pojkar klättrar på trästolpar i en smutsig flod.
En äldre afroamerikansk man i gul skjorta står framför ett informationsställ.
Tre äldre kvinnor går bakifrån.
En man med ögonbindel siktar på en pinata medan folk tittar från däcket bakom honom.
Man i orange skjorta hukar och arbetar på svart cykel.
En kvinna i svart klänning står bredvid en rosa cykel.
Mannen i vitt städar golvet.
En kvinna målar en bild av en stor byggnad som syns i bakgrunden.
Barn läser och skriver.
En man med ryggsäck och en promenadstav utforskar en bergig terräng.
Män arbetar på en byggarbetsplats.
En grupp kvinnor, som ser olyckliga ut, sitter i ett kök och pratar.
Två personer sitter på en klippa med utsikt över floden.
En man sitter på gräset och håller ett barn framför sig.
En man sågar genom en träbit för att reparera ett stängsel.
Band som spelar framför en liten publik utanför.
En liten pojke som leker med ett hjul.
Två unga svarta män i blå jeans sitter framför en hängmatta.
En grupp människor går nerför en lantgata.
Två asiatiska kvinnor utför uppgifter och det finns en vacker bakgrund av bambu.
Tre stora hundar springer snabbt bredvid ett hus.
En grupp kvinnor går nerför gatan med öppna paraplyer för att skydda dem från regnet som kommer ner från himlen.
Kvinna som gör sushi på köksdisken.
Den bruna hunden går genom en flod omgiven av buskar.
En ung afrikansk flicka i en vit stol gör en annan flickas hår.
Ett afrikanskt amerikanskt barn i röd flanellskjorta sover på en vävd hängmatta.
En liten pojke glider ner för en röd rutschkana.
En kvinna i grön klänning som röker en cigarett dansar med en partner.
Två unga män hoppar över två stora trästockar.
En man som sätter en liten pojke i orange i en barngunga.
Två män slåss när de spelar frisbee.
En leende kvinna i en orange kjol har en öppen portfölj som visar en klohammare.
En kille som instruerar folk bakom tåget.
En man i grön skjorta håller en böljande nål medan han röker en cigarett i ett rörigt kök.
En man som använder en kran koncentrerar sig i en skyddande monter.
Två personer sitter i en lång träbåt i en vattensamling.
Ett ungt par njuter av några snökoner på trånga gatan.
En ung man kastar upp en svetsarmask när en ung flicka tittar på, en sex-pack, grill och krita meddelande i bakgrunden.
Folk står på en tågplattform och väntar på tåget.
En sovande bebis i en haklapp som ligger på en filt.
En svart man, på en trottoar, spelar dragspel.
En man sitter vid ett bord och äter och dricker.
Två dykare interagerar med en delfin under vattnet.
Tre kvinnor utanför alla klär sig likadant och pratar med varandra.
Svarta kvinnor gör tyger i sitt hem.
En man med medellångt hår, bär en röd mössa och blå shorts utan skjorta, på ett knä på stranden, skulptera ett sandslott med en tråg.
Blond pojke äter en smörgås på en vit stol.
Ett gäng cowboys väntar på sin utmaning att fånga ett levande djur.
En grupp människor i vitt stånd med vita getter.
En man och en kvinna delar en kyss på stranden.
Kvinnan städar fönster framför butiken.
Gatudans på plast medan en stor grupp ungdomar står och tittar på.
En quarterback är på väg att kasta ett pass från slutzonen i en fotbollsmatch.
En liten flicka kramar sin bror på en gångbro i en skog.
En flicka går utför förbi några parkerade bilar.
En pojke försöker sätta en skärm på ett fönster.
En ung svart man med två vapen riktade mot huvudet.
En kvartsback, i frihetsstatyn, hålls fast av en motståndare bakifrån.
Hunden jagar geten runt gården.
Man i rak jacka försöker komma loss, står framför barn med Jenga block.
Pojken är i poolen med en vuxen kvinna.
En glest befolkad arkad med många ljust upplysta spel och några personer strödda runt.
En man som bär kamouflage styr en motorcykel över några stenar.
Fyra unga män njuter av ett dopp i den lokala sjön.
En familj sitter i en park på gräset.
Ett pepband i röd och vit uniform spelar när man sitter på en stadion.
Kvinna med rött lockigt hår tar bilder utanför.
En kvinna som rider en häst på en jordarena, bär på en amerikansk flagga.
En liten flicka visar sin bror tillgivenhet.
Tre unga flickor klädda i vita klänningar springer mot en fontän.
En kvinna och ett barn som går förbi en vandaliserad byggnad.
En ung flicka och en hund bredvid henne tittar på något i en bäck.
En liten flicka kastar stenar i en bäck.
En mycket ung blond tjej med rosa byxor med vita prickar sitter på en skogsstig i en skog.
Hunden står i vattnet bredvid gräset.
En man i en blå långärmad jacka som skriker av rädsla.
En kvinna med shoppingväskor går förbi tunnelbanan.
En flicka i rutig klänning går på en trottoar bredvid en stenbyggnad.
En grupp i kostym sjunger på en renässansmässa.
Två kvinnor spelar tangentbord under ett upplyst tält på natten.
Folk på ett betongområde tar bilder.
En liten pojke ler och pekar medan en man tittar i barnets blickriktning.
Den bruna hunden är på väg att bita en tass tryckt boll.
Två män i svarta skjortor som står på ena armen.
Bakverkskockar är på väg att sortera bakverk.
En man klädd i rött och vitt spelar banjo medan andra ser på.
En grupp leende unga kvinnor poserar tillsammans.
En kvinna med mörkt hår håller en grönsak när hon står framför ett bord fullt av grönsaker.
En man och en kvinna dansar på gatan.
En man håller i ett utensil och gör sig redo att gräva i en tallrik fylld med mat.
Två hundar brottas i marken.
Fyra män åker rullskridskor i en kö, och de tre sista håller i höfterna på mannen framför dem.
En kvinna på en mörk bar som pratar med folk.
En ung blond tjej i rosa skjorta och grissvans sitter ovanpå en mans axlar i en publik.
Mannen hänger upp en bild av trädet när kvinnan tittar på.
Två barn leker och en man i svart byxa går nära barn.
En mager hund springer genom grönt gräs.
Tre mellanöstra män i affärskläder sitter runt ett bord.
En flicka i rosa snurrar ett band.
En blond kvinna erbjuder ett fat mat till en annan blond kvinna medan hon sitter vid ett vitt bord.
Man tittar in i kameran och spelar gitarr
En gammal man i arméutmattning riktar uppmärksamheten på en rad barn som står i fokus.
En flicka hoppar i gräset.
En man i grön skjorta skrattar bredvid en kvinna i gul tröja, håller i en rosa ballong och bär en rosa tiara.
Tre hundar springer ner i vattnet.
Två unga flickor springer över ett fält när de flyger en drake i den molntäckta himlen.
En arbetare som ser till att hans maskin fungerar korrekt.
En man som bär en grön jacka svetsar en stor metallbit.
En svetsare i masksvetsning med gnistor som flyger.
En liten pojke med svart lockigt hår sitter i en blå stol som är på trottoaren.
Gråvit man med glasögon, använder smed verktyg.
En ung pojke i röd skjorta pekar på något.
En grupp på 4 personer arbetar med mycket papper.
En ung man är i en bäck med sin smutscykel.
Fyra män tittar på ett stort tecken.
Tre män på en ställning som uppförts utanför en byggnad.
En lerig gyllene hund som springer i gräs
Två barn springer i sanden, längs stranden.
En hund springer med en gul tennisboll och bär en röd sele.
En man som bara har underkläder och tennisskor på gatan.
En svart hund springer genom vattnet.
En liten hund hoppar i vattnet.
Tre unga pojkar hoppar och leker i höet.
En man håller metallfälgar en med varje hand medan han pratar med två personer.
En ung man med bruna ögon är klädd som Jack Sparrow.
En man med en tanktopp som håller upp en skylt som introducerar Mark Finley.
En ung pojke glider på gräset i ett innerrör
En brun fågel sitter på en trädgren.
En man i gul skjorta klädd i mångfärgade plastsmycken.
En man i morgonrock rider en åsna nerför en gata.
En man håller en bok framför en krittavla.
En ung flicka och en äldre gentleman håller hand när han pekar på något utanför ramen.
Männen pratar med personen i polisbilen.
En konstnär som arbetar hårt för att rita ett komiskt porträtt.
Ett gammalt par går upp för en sandhög.
En person hjälper en annan person upp till toppen av en sandhög under en molnig himmel.
Två fordon står parkerade utanför en liten livsmedelsbutik.
Variation är livets krydda oavsett vad kulturen kan vara.
En buss som en mekaniker jobbar på.
En arbetare som står på en hög ställning.
Män utför vägarbete mot en bakgrund av bruna kullar.
En man i en blå kanotpaddling i havet.
En del människor står ensamma på stranden i sina baddräkter.
En man i svart skjorta och röda shorts sitter på stranden av en sjö.
En lärare som visar sina elever något på en projektorskärm.
En kvinna och en ung flicka hänger kläder på linjen.
Två vandrare vilar på ett snötäckt berg.
En mycket stor grupp människor står utomhus under de vackra molnen.
Person som läser ur en bok för ett rum fullt av människor.
En man sitter på en bro vid en flod och spelar dragspel.
En del byggnadsarbetare är på en plattform och arbetar till en byggnad.
En brevbärare i sin lastbil som står framför en grind.
Ett barn som sover i en bil med fönstret öppet
En ung flicka med lockigt hår med vit skjorta med skalle och benbild på.
En ung flicka gör ett fånigt ansikte för kameran.
En man som bär orange skyddsväst och en hatt använder byggutrustning.
Pojke med röd jacka gör ett handstånd på gräset.
Ett litet barn springer mot kameran i en park.
En hund och en dammstorm.
En äldre kvinna med en näsduk och en käpp står på en slaskig kullerstensgata.
En man med ett leende som sitter på golvet och lagar sin cykel.
En grupp människor står och samtalar inne i en byggnad.
En man står på röd ställning.
En man med arbetshandskar och verktygsbälte klättrar uppför ställningen bredvid en gammal gul och vit byggnad.
Två barn tittar på något spännande som en vuxen visar dem.
Två män försöker skrapa cementen från golvet för att jämna den.
Ett band som spelar på en gata som åskådare klocka
En skateboardare klädd i svarta jeans, vit t-shirt och röd bollmössa kommer från läppen på en ramp och suspenderas i luften.
Fyra personer framför Wells Fargo.
Två personer håller ihop sina händer över en tredjedel, framför en upplyst scen.
Ett barn, som bär grönt, studsar på studsmattan.
En grupp collegestudenter samlas i communitycentret.
En familj vandrar över ett stenigt landskap.
En grupp fans på en stadion bär rött och hejar.
En kvinna som njuter av att läsa på ett kafé
En afroamerikansk man tittar genom ett mikroskop och det finns en affisch där det står blodceller hängande på väggen.
Tre personer leker i snötäckta stadsgator.
Två pojkar sparkar en boll mot varandra i parken.
Män klädda i drag utanför en affär.
En pojke lägger sig med en orange boll framför en rad blå bilar.
Ett kvinnligt barn med en handduk bredvid ett handfat.
En kvinna borstar bort damm och smuts från ett möjligt fynd.
En hund springer på ett fält.
Toddler sitter i en gunga vid parken med en gul sippy kopp.
Ett par pratar med en man som sitter med en hammare.
Två paraglidare övar sin farkost på ett öppet fält.
Ett barn med cowboyhatt som springer mot ett annat barn.
En ung pojke försöker plocka upp en pumpa i en pumpaplåster.
Folk i asiatisk dräkt går i en parad.
En mager brun hund går över ett stort stycke fallet träd.
En man som jobbar på ett fönster i den gamla byggnaden.
En man tittar in i spegeln och rakar sig medan en kvinna tar en bild av honom.
En pojke är märkligt uppmärksam på skor.
En man med blå skjorta, blå hatt och förkläde står utanför Candy Cafe en solig dag.
En flicka sitter på stranden och stirrar på havet.
Den bruna och vita hunden niperar mot den gula hunden.
Flicka med solglasögon och shoppare i en liten affär.
En man med en konstig hjälm sitter ovanpå en blå motorcykel.
Ett litet barn sover medan det håller ett uppstoppat djur.
En äldre man som sitter emot ett samtal med en gitarr i sina händer.
Det finns tre personer som bär dräkter, av vilka två spelar blåsinstrument.
En man spelar fiol utanför på en trottoar.
En man, i en svart tröja, fiskar.
En man som reparerar ett cykeldäck medan hans kund ställer frågor till honom.
En publik står på gatan.
Föräldrar som lär ett litet barn att åka skridskor.
En ung pojke hoppar ner för en uppblåsbar vattentur.
En ung pojke som står på en gunga framför en blå rutschkana.
Daredevils njuter av bergsstigning nerför ravinen.
Två äldre män, i ett vitt rum, leker med en marmorskulptur.
En liten flicka i en swing skrattar.
Ett band bestående av två män och en kvinna spelar för en grupp människor.
Två män med rakade huvuden, båda bär vita skjortor utövar undervattensdykning.
Två konkurrenter, varav en i USA:s flygvapen, brottas.
Några barn i barnvagn undrar mycket.
Två män hanterar en grå hund med ett blått knutet rep i munnen.
Man sparkar fotboll av tee i t-shirt och shorts
En man med kanot är på stranden med tält uppsatt.
En skjortlös man som lagar mat medan han campar på stranden.
En del joggar ute i mörkret.
En liten flicka leker i höet.
En man somnade när han läste Da Vinci-koden.
En man med blå byxor böjer sig över för att plocka upp något från marken
En man i Alaskas tröja och keps köper lotter.
Två män bygger något tillsammans.
En flicka leker med ett halsband när solen skiner bakom henne.
En liten vit hund tigger.
En liten flicka som sitter på golvet och håller i gitarrhandtag.
En man i glas grillar korv och köttbiffar på en grill.
En pojke i röd hatt tar bilder med sin kamera.
Ett litet barn som tar en bild med en kamera på ett stativ.
En kvinna i vit skjorta och rosa byxor står bakom ett bord med tårta, jordgubbar och slag.
En kvinna som öppnar en present runt sina vänner.
Två grå hundar och en svart hund som leker i en damm under en överfart.
Det sitter en kvinna vid ett bord vid köket.
Tre personer på ett tåg som håller spelkort, ler.
Två hundar och en valp.
En man sprutar en vätska från en lång slang på stranden.
Flera personer gör en synkroniserad dans med hoppning.
En liten pojke placerar föremål från en vagn på kassan.
En man klädd i en glänsande astronautdräkt poserar för en fotograf på en trottoar.
En ung man i blå skjorta har armen runt en ung kvinna i en röd jacka.
En flicka klättrar på ett djungelgym.
Asiatiska barn klädda i rött och gult, och bär svarta knäskydd, rullskridskor utomhus över stora, glänsande kakel.
Tre pojkar spelar tagg på stranden.
En flicka med upplyfta armar glider nerför en röd och vit rutschkana.
Tre simmare simmar eller tävlar i separata körfält.
En stor grupp människor i röda soldatjackor står i kö utanför.
En pojke hoppar från toppen av ett blått plastglas.
En man i rutiga byxor svart jacka och en rutig hatt håller en servitör bricka.
En bergsklättrare i en röd hjälm tittar nerför klippan.
En kille i en hård hatt som jobbar på några maskiner.
En kille som pekar på en jättestor björnbär.
En grupp kvinnor som går med väskor på axlarna.
En man och en kvinna är utanför en bil som är fylld med föremål.
En ung pojke och flicka som spelar baseball på ett gräsfält.
En stor publik leker i och runt en fontän.
Bilden är av ett centrum område med människor korsar gatan, och promenader på trottoaren.
En kvinna i sweatpants står vid toaletterna.
En kvinna och hennes dotter mäter sig mot en jättehärskare på "Washington Farms".
Flera män, alla klädda i rött, drar på sig ett rep.
En grupp människor som sitter på betongtrappor på en basketplan i grannskapet.
En blond tjej som öppnar ett grönt paket.
Man i en topp hatt, spelar sitt dragspel på trottoaren vid en gata
En kvinna som uppträder genom att sjunga en sång.
En skallig man med en blå skjorta som äter revben vid ett bord utanför.
Mannen står på kanten av stor klippa med utsikt över naturskön utsikt.
En man läser upp ett pappersark för en folkmassa medan en annan man i vitt står bredvid honom.
Pojke i bubbelbad, skrikande eller sjungande till skrubbborste.
En grupp ungdomar sitter utanför och lyssnar på en gitarr och fiol som spelas.
En ung pojke kryper med ett litet barn.
En man bär ett förkläde som står i köket och håller en tallrik.
En pojke håller upp en röd hink till en ponny.
Preteen flicka med blont hår leker med bubblor nära en försäljare stall på en köpcentrum gårdsplan.
En kille i kostym som leker säckpipa bredvid en tjej som bär tölplagg.
En hund försöker fånga en snöboll i munnen.
Du måste svara din chef.
En person som sätter upp ett tält bredvid några andra tält på den snöiga marken.
Ett par som håller händer stannar för att titta på något.
En ung pojke leker på en lekplats bit formad som en sjöhäst.
En ung pojke simmar i en pool.
En pojke utan tröja och volleyboll i handen.
En grupp skolbarn går upp på en lantväg på hösten.
Ett kvinnligt barn sprider Nesquik pulver på ett bord.
En man i cowboystövlar, kalsonger och gitarr håller i en kvinnas arm.
En ung asiatisk man som studerar med en penna och en ordbok medan han dricker en cola.
Få människor liftar på baksidan av en sopbil.
En man är en grön skjorta rör om en skål med mix nära en spis med två stekpannor.
Flera unga kvinnor går längs en vacker korridor
Två asiatiska kvinnor och en ung asiatisk flicka med trehjuling står utanför i skuggan.
En liten pojke som försöker klättra upp.
En ung pojke i en blå jacka drar upp något svart ur en tygpåse.
En pojke lagar hjulet på sin cykel.
En man med blå skjorta och röd hatt ridande på baksidan av en vagn fylld med hö och dragen av en vit häst.
Fem män på en restaurang poserar för en bild.
Två kvinnor i vita klänningar går förbi en annons med två golfare på den.
En kvinna går vid en flod över stadsbyggnader.
En spelare på det vita och blå laget sparkar en fotboll mot sin lagkamrat medan spelare på det röda laget klocka.
En hund hoppar på damen medan den andra går sin väg.
En hund vilar i ett gräsfält
Killen rider en stor brun tjur.
En asiatisk kvinna i gul skjorta tittar på vykort medan hon är i kassan.
En brun hund som leker i lera.
Massor av människor som spelar en vatten shooter karneval spel.
Två personer bär hjälmar som har ljus på toppen.
En flicka med svart hår och tandställning bär solglasögon och poserar med en trärobot.
En kvinna som sitter i en tvättomat och tittar på kameran.
En person med en mängd olika varor som står bland flera andra på en grusväg.
En man som går med ett badkar av något på huvudet.
Flera personer går upp och ner för en trappa i en gränd med graffiti målad på väggarna
Publiken njuter av stranden.
En man i en basebollkeps spelar ett skjutspel i en arkad med en vän.
En grupp människor gör ett projekt för en frivillig organisation.
Två fotbollsspelare blir insnärjda medan de båda går för bollen.
En ung man som skateboardar framför havet.
En kvinna med en svart skjorta som pratar på sin mobil när hon går på en väg.
En svart kvinna går mot en kvinna med gul hatt.
Musikern i den bruna rocken går i sina tennisskor.
En kvinna som bär antikviteter, däribland många pärlor.
Ett par sitter på motorhuven i en bil med ryggen mot kameran.
En bil är delvis nedsänkt i en sjö.
Tre kvinnor som bär svart är bredvid varandra på ett tåg.
En man sitter på en segelbåt och solen går ner bakom honom.
En liten pojke undersöker ett par blå jeans, med en vuxen i bakgrunden.
Scenen av en olycka där en buss körde på en mc.
En liten flicka i röd klänning står på en stig i skogen med en häst i bakgrunden.
Folk i kostym står runt ett träd i en skog.
En ung flicka springer på en strand bakom en ung kvinna som sitter och spelar gitarr.
En kvinna som ger ett litet barn en röd skjorta ett föremål från en inköpskorg.
En byggnadsarbetare håller upp en stoppskylt för att flagga ner trafiken.
En man jobbar i en affär med munkar.
En mans händer håller en bit metall på ett sliphjul.
Blond kvinna som röker en cigarett i sina väskor.
Två män med verktygsbälten sätter fast en skylt i en byggnad.
Två personer poserar för kameran.
Grupp av personer som sitter vid röd stol och bord.
En grupp människor protesterar genom att sälja människor.
Två män trycker på en lastbil som har en bild på en kvinna på sig.
En man står på sin kolgrill.
En man i hatt med grön skoter står vid vattnet i en park.
En motorcykelförare svänger till vänster.
En kvinna lutar sig mot stolen och spelar elgitarr.
En man sjunger medan en annan spelar gitarr under en scenföreställning.
En man håller en gitarr på en livlig gata medan folk tittar på.
Kvinnan sjunger på en klubb under starkt ljus
En kvinna i blå skjorta och svarta byxor går längs en väg.
Två gatukonstnärer uppträder på trappan för en grupp åskådare.
En kör står upp på ett podi som sjunger en sång.
Folk skriver under i en kyrka.
En blandad könskör i mellanstorlek sjunger medan regissören motionerar för att hålla takten.
En fläckig hund hoppar över en lerig bäck.
En arbetare som bär en ljus väst och svarta kläder plockar upp sopor på marken medan folk går över gatan bakom honom.
En flicka på en strand med regnbågsflaggor.
En man i en simbassäng håller en leende pojke i en flytapparat.
Det här är baby, klädd i blått, stående barfota på en sten.
En unge med gröna skor, röda shorts och en blå hatt och skjorta står på en sträcka av trottoaren.
En brun hund som travar över en gräsbevuxen inhägnad gård.
En liten flicka sitter ovanpå en pumpa framför ett arrangemang av levande blommor utanför.
Fyra soldater går och pratar med varandra medan de håller i vapen.
Två män i vandringsstövlar slår kampsporter poser.
En kvinna och en man njuter av sin drink på festkvällen.
En äldre man med en "slow" skylt ler mot kameran.
En hund som ska hoppa för att fånga en frisbee
En brun hund hoppar upp i luften för att fånga en boll.
Tjejen slår en fotbollsboll under en match.
Två män delar ett samtal mitt i en park, bakom ett kort staket.
Två män i svarta skjortor samtalar runt en videokamera.
Två män arbetar tillsammans för att intervjua en sittande man på en stor teater.
Folk håller skyltar och marscherar.
En kvinna på scenen som håller en mikrofon stående av en man.
Två asiatiska män ler samtidigt som de firar en födelsedag med en lager chokladkaka med ett gnistrande ljus.
En man i en grön hatt är böjd över sin DJ-utrustning plugga i en mikrofon
En man håller en stående kvinnas fot med båda händerna.
Tre kvinnor i zigenarkjolar står runt parkeringsplatsen för Notre Dame i Frankrike.
En kvinna som skrattar i en bar.
En liten gata med några personer som går nerför den.
Två barn vid ett träd nära lite vatten.
En flicka i rosa står framför en Mud kaffebil.
Detta är bilden av två asiatiska män som hukar sig nära en mopp-pad.
Fotgängare och bilar tar sig genom Times Square i New York.
En man hjälper ett litet barn att komma på ett tåg.
Tre sittande människor äter och dricker nära träd, och tre personer står i bakgrunden.
En man som står framför en grind inne i en kulle.
En man och en kvinna som dricker och roar sig på en nattklubb i staden Angeles.
Tre barn sitter runt ett bord och läser böcker.
En pojke står bredvid en bil framför en klädstreck.
Folk sitter i en hörsal med program.
Två kvinnor böjde sig ner och arbetade ute på fältet med träd i bakgrunden.
Mycket många skidåkare är samlade på en skidplats.
Folk går genom ett snötäckt fält med ett berg i bakgrunden.
En vuxen hjälper ett litet barn att laga sina glasögon.
En kvinna med vitt visir och blå topp och vita byxor som äter medan hon står i folkmassan.
Ung pojke i baseballuniform knäböjer för att fånga en boll på ett baseballfält.
En man med långt hår och en blå skjorta sitter ute med sitt gitarrfodral öppet och skrattar när en ung flicka sitter och tittar.
En kvinna bär en korg på huvudet bort från vattnet.
En hund sniffar en nyskuren trädstam.
Två hundar leker i gräset.
Etniska människor besöker plocka färsk mat att köpa.
En kvinna springer på stranden.
Tre kvinnor, klädda för ett formellt tillfälle, tar sig en stund att le.
En hund som hoppar genom en svart och vit båge.
En man som säljer färgstarkt mönstrade mattor njuter av en drink från en kaffekopp en solig dag.
En man med långt mörkt hår och mustasch går nerför gatan i shorts och cowboyhatt.
En motorcykelförare klädd i orange växel svänger till höger.
En man bär ett tecken medan han står i regnet.
En man skalar ett rent rockansikte med repstöd.
Fyra campare njuter av en kväll runt en vedeld.
En motorcyklist med en röd hjälm kör sin blå motorcykel nerför vägen.
Tre män går utanför en vit byggnad.
Två orientaliska ödlor kämpar för dominans i en liten damm
Människan använder uppblåsbara leksak för att spela en gräsmatta spel.
En grupp rasbuggies färdas längs en kapplöpningsbana.
En person med tatueringar på armen med motorcykelhjälm.
En familj och vänner sitter och äter vid ett bord fyllt med många skålar med god mat.
En collie springer nerför en rutschbana.
En man med brun jacka står bland en grupp män framför en stor maskin.
Folk som klättrar i trappor till en plattform.
Två män i en bar gör lustiga ansikten medan de håller en drink med sin högra hand.
En skallig man i vit skjorta dricker ett glas öl.
Mannen i en blå skjorta, med hjälm, är redo att klättra.
En man som borrar hål i en pumpa.
En man filmar en annan man som börjar klättra upp för en metallstruktur.
En man som förbereder sig för att stöta bort ett berg.
En medelålders kvinna klädd i en röd kjol, brun blus engagerad i att göra keramik.
En man står nära ett kristet tecken, när ett offentligt tåg passerar bakom honom.
En hund hoppar och fångar en frisbee i gräset.
Unga vuxna har grillfest i parken.
En man med vit jacka håller i en svart bok.
En man som fiskar från stranden på vintern.
En man och en kvinna tittar på utsikten på en trappa vid havet.
Baby med orange skjorta och matchande pannband med ett brett leende.
En ung vit man med kort skägg rockar ut på sin gitarr.
En kvinna som rörde vid en mans ansikte på en vägg efter att de tagit en paus från att köra motorcyklar.
En vuxen kvinna och ett ungt gossebarn som går längs en pir och håller i ett paraply medan det regnar.
En skolpojke, med ryggsäck på, hoppar från en vägg.
En leende man i vit skjorta grillar på en öppen grill.
En vit hund som tittar på en svart hund i luften.
En svart hund hoppar för att fånga en boll i munnen nära en stenvägg.
En man som läser en tidning i ett tåg.
En hund som ligger ner, fastbunden vid sidospegeln på en gul VW-buss.
Två män sitter på en bänk mellan två träd med utsikt över ett höstlandskap.
Pojken träffar den blå och vita fotbollen med knäet.
En man observerar uppmärksamt en bild genom ett mikroskop.
Ett barn tittar upp på en vuxen medan det sitter i en barnvagn på en trottoar i staden.
En liten flicka i en gunga skrattar.
En grupp på sju personer äter vid ett bord som är garderat i en svart duk.
Två män hugger ner ogräs på gården.
En man i röd rock kör ett fordon.
Kvinna och liten svart hund går över trottoaren
En grupp barn springer i gräset.
En man i lila, vitt och gult på styltor.
En man i söndersliten skjorta och byxor, sitter på en stol och väver något.
Mannen i blommig kostym och hatt uppträder med hula-hoop i staden gatan.
En man som bär grön jacka och stickad hatt sorterar tomater på en utomhusmarknad.
Två hundar springer genom surfingen.
En hund springer genom högt gräs med en kvinna klädd i rött i bakgrunden.
En kvinna som väntar på nåt på trottoaren.
En man sitter på trottoaren framför en asiatisk restaurang när folk passerar.
En grupp människor som stod runt två män sittandes i turbaner.
En målvakt försöker blockera en puck hit av en spelare på en ishockey spel.
En asiatisk kvinna cyklar framför två bilar.
En kvinna som sitter vid ett bord stickar och tittar på en hockeymatch på TV.
En kvinna arbetar ett projekt med tråd i handen.
En pojke försöker kyssa en annan i ett skollunchrum.
Passagerarna på bussen är uttråkade.
En äldre man som bär hatt och jacka cyklar nerför en stenlagd stig medan solljuset strömmar genom höstträden framåt.
En grupp människor som arbetar vid ett konferensbord, på ett kontor.
Asiatisk man i kostym och glasögon tar en tupplur vid dörrarna i en tunnelbana.
En pojke tittar ner och breder ut sina armar
En grupp människor klädda i blå skjortor, stående i gräset.
En bicyklist och en man i kostym sitter nära en fontän och pratar på mobiler.
En vacker långhårig blond tjej klädd i en blå och grön bikini som går nerför en gata
En gatuartist med vitt ansikte ser folk gå förbi.
En rad människor som går genom en torr region förbi en skylt, människor antingen går eller rider djur.
Ett gift par sitter i ett fordon.
Flera motorcyklar är parkerade på en parkeringsplats.
En liten flicka glider ner för en spiralbild på lekplatsen.
Två män som jobbar utomhus och städar gatan i sina orange uniformer.
En polis visas arbeta en blockparty.
En hane står på en bas och kastar en boll.
Två unga flickor rider röda trehjulingar.
En vacker kvinna som dansar på en parad som håller i en liten pojke.
Många klädda i arméutrustning går på kraschen går en brun hund.
En man i en militäruniform står bredvid vad som verkar vara en militär k-9 hund, med en högtalare i förgrunden, och annan militär personal och militära fordon i bakgrunden.
Man tar en bild i en skara människor.
En man och en kvinna går genom gatan under en parad.
En grupp människor tävlar i loppet om ett botemedel.
En stor grupp människor går för en sak.
En fiskare arbetar på nätet medan han är på land.
En grupp människor rider på en John Deere traktor på ett fält.
Det finns en grupp små barn några bär ryggsäckar sitter på en kulle.
En grupp människor rider på ett tåg medan de tittar ut genom ett fönster.
En man och ett barn som poserar framför ett tåg.
Den lilla pojken i den röda skjortan stack huvudet ut genom fönstret på tåget.
Folk går på en trottoar förbi ett parkerat tåg.
Små barn och vuxna går runt plattform 9 bredvid tåget.
Tre kvinnor chattar medan de sitter i ett väntrum.
En kvinna i rosa jacka går förbi ett skyltfönster med en röd klänning i en urban miljö.
En person som läser något sitter under trädet.
2 män målar en träbänk utanför.
Två sköterskor som sitter på en bänk och väntar på en buss.
En man står bredvid en röd dörr.
En äldre arbetare står i våt cement med en tramp.
En man i blå skjorta står i en dörröppning.
En man som håller en kamera under vattnet.
En brun hund möter en svart hund och en vit hund på ett fält av långt gräs.
Tre hundar springer genom ett gräsfält.
Många människor står på en buss med ljusa gula overhead handtag.
En liten pojke skakar snön av ett träd.
Ett yngre barn som bär en röd tröja som visar vad han har i handen.
En man som borrar hål i en metallbehållare.
En hund som går längs en sprucken och ashen yta.
Sju personer sitter runt ett svart bord och spelar kortspel.
En man i svart skjorta och glasögon skär en tomat vid ett köksbord.
Unga pojkar tar hem lite frukt.
Crouching Man i alla vita skjorta och byxor arbetar med en stor vävstol.
En man som plockar upp en stor sten.
Två personer i forsränningsredskap står på en torr, stenig flodbank, som pekar mot floden.
En pojke sparkar en boll när andra barn tittar på honom.
Fyra äldre kvinnor sitter och talar på en parkbänk.
Mannen i vit skjorta och bruna byxor sätter nya bältros på taket.
Byggarbetare i gult och orange arbete på en stad gata.
En man trycker ner ett fyrhjuligt kort på gatan.
En man som bär en röd livväst vågor som han vattenskidor.
Person i röd skidjacka skidåkning baklänges
En man som bär en röd flytväst åker vattenskidor över en vik.
Ett barn med och vuxen hand.
En flicka står bredvid en cykel parkerad framför en byggnad medan två män, en med gitarr, går förbi.
Två unga pojkar som spelar schack i ett rum.
Människor i en hamn tar emot och fraktar ut varor nära en trevlig stor vit båt.
En kvinna sitter i klippor vid havet.
En fiskare fiskar vid stranden av en dimmig flod.
En man spelar gitarr på stranden.
I detta förvrängda foto visas en man på en grusväg med en hopphund.
Ung man skalar citron med en kniv i en röd korg.
En svart hund hoppar upp ur vattnet.
Grupp av deltagare går bakom flyt i asiatiska parad.
Två människor som sitter med dreadlocks.
En byggnadsarbetare byggnad väggar med en borr.
Ett par står högst upp i trappan och två personer står längst ner.
Musikkonserten har precis startat på Giant stadion
Trafikpolisen styr trafiken framför en bil med ohio-plattor på sig.
En blond man sjunger passionerat in i mikrofonen.
En person med en flerfärgad hatt står precis bakom en mosaik med spanska ord och framför en gräsbevuxen kulle.
Två kvinnor flyter i en Busch Gardens fat genom en slingrande vattentur.
En kvinnlig cyklist klädd i rött använder en kommunikationsapparat medan en annan går förbi.
Två män väntar i gathörnet trots att det regnar.
Två män i svarta rockar står vid sidan av en byggnad.
En man i röd skjorta spelar elgitarr.
En grupp vuxna och barn befinner sig på en nöjespark och vakar över ett räcke.
En man knuffar ett barn på ett leksakståg.
Bum lyssnar på radion vid en ljus stolpe nära stranden.
En liten flicka går in i en pool.
En pojke och en medelålders kvinna går ut från en folkmassa utanför.
En man och en pojke smakar frukt.
En man och en kvinna njuter av en trevlig måltid på en utomhusrestaurang.
En man i gul skjorta sågar plywood.
En kvinna i blå, solbränd och beige randig skjorta röker.
En ung man står i köket och håller i en stor gryta.
En man i röd skjorta och en kvinna i en färgglad skjorta och sitter utanför.
En livlig karateträning på dojo.
Ett ungt barn som bär grönt leker med vakuumslangen på golvet.
En man och en kvinna diskar i ett kök.
En vit manlig underhållare på gatan bär en svart skjorta och blå hatt med en gul rand.
En konstnär som målar väggen täckt av bambu.
Mannen i svart skjorta kramande kvinna i vit skjorta, grå kjol.
En flicka med rosa skjorta springer genom blommigt gräs.
Några turister tar bilder på sina hundar med den molniga himlen som bakgrund.
En man som spelar gitarr och sjunger utomhus.
En man i blå skjorta och en kvinna i klänning som har ett samtal medan han dricker.
Två personer bär en korg fylld med mat nerför gränden.
Medan man sitter på en stol, blåser en man i en blå skjorta, grå byxor, mångfärgade bandanna och inga skor genom ett långt rör.
Byggarbetare som fixar järnvägsspåret.
En byggnadsarbetare gör en del slipning på en bit järn.
Två kvinnor som leker och ler.
Arbetare i reflekterande kläder med spadar på tågspår.
Två kvinnor går förbi en affär och tittar in.
En mor står i ett kök och håller ett litet barn.
En ung pojke sitter på gräset.
Två män pratar om affärer över öl.
Två kvinnor med brunt hår prat.
En kvinna som bär en babushka sitter och sover inne i en blomsteraffär.
En grupp människor arbetar på en sandskulptur.
Det finns en grupp människor och en svart hund i ett vardagsrum och matsal, några sover lite äta.
Fysiskt utmanad person som sitter på sin rullstol i en park.
Ett barn sover på en soffa med munnen öppen och handen draperad över bröstet.
Fem vuxna sitter på stentrappor.
En ung kvinna i en grön blus med en plastpåse stående på tunnelbanan.
Butiken var öppen trots att en man arbetade på byggnaden.
En man på jobbet gör ett litet svetsjobb med ett lödverktyg.
En brun och vit hund travar längs vägen på hösten.
En ung person med en mohawk och en näsa piercing i en rutig skjorta.
En man i lila jacka har ett uttryck i ansiktet.
En äldre kvinna som bär baddräkt håller en picketskylt medan hon deltar i en demonstration om invandring.
En bongospelare med röd skjorta som spelar i ett band.
Två fotbollslag på en fotbollsplan med domaren.
Tre pojkar som spelar fotboll.
Två pojkar står mitt på gatan, den med svarta shorts står och klappar ihop händerna medan den andra i grått springer framåt.
En pojke springer på trottoaren framför en blå byggnad.
En svart och vit hund leker i vattnet.
Ett barn på en falsk hästtur.
En man med mikrofon läser ur ett papper när han står framför två män som håller i tubas.
En publik ser en hund klättra uppför en trappa.
En kvinna sitter på en grå bänk framför en betongvägg med graffiti.
En man som bär svart skjorta och jeans bowlar med boll och 9 sprayburkar.
En kvinna i mörkblå T-shirt väver ett randigt material.
En antilop löper genom högt brunt gräs.
En dam som bär bollmössa lär sig att väva tyg av en kvinnlig instruktör.
En gatuartist med gitarr.
Två män bär svarta västar och vita skjortor och en flicka håller flaskor med öl.
Två personer sammanflätade längs en cementgång.
Två flickor går längs gatan och pratar.
Mannen i kostym tar en tupplur i parken.
En liten pojke med blå balans när han går på en stor klippa.
Två hundar leker på gräs.
Tre män sitter utanför framför en byggnad, och var och en spelar ett instrument.
Cheerleaders är på fältet och hejar på.
Mexikanska kvinnor i dekorativa vita klänningar utför en dans som en del av en parad.
Två män med rockar och vapen som bär en död kanin.
En man i kostym står på gatan med sin högra hand utsträckt.
Mannen vinkar till sin familj från toppen av bron.
Bilden är av en kvinna som tävlar i ett lopp som gör backstroke.
Tre män njuter av ett gott skratt.
Två män i ljusa skjortor och mörka byxor sitter på en balkong och samtalar när en ensam bil passerar nedanför.
En kvinna i rosa bikini bredvid en man i brunt.
En kvinna som går i bikini mot en man i randig skjorta.
Kunderna står i kö vid en maträtt.
Damen ber hunden att ge henne bollen på deras strandpromenad.
Två barn i en leksaksbil på en bensinstation.
Tre barn leker på en grusväg i naturen.
En kvinna som väntar vid tågspåren.
Två damer går över en gata framför en restaurang.
En kille paddlar genom några forsar.
En man i vit skjorta och svarta byxor står med vänster hand på huvudet.
Asiatiska barn som leker med en rail.
3 barn med hattar som leker på en häst
En liten flicka poserar på sin cykel med sin hund i skogen.
Ett litet barn som kramas av en kvinna med ljusbrunt hår.
Män med säckpipa och kilt står runt i en cirkel.
Tre män i kamouflagekläder och en annan man i hatt och röd skjorta och blå shorts står framför en byggnad.
Mannen i randig skjorta tar en bild av den andra mannen i grått.
Två gamla män sitter bredvid en ung asiatisk kvinna i konstiga stolar.
Barn klädda i Halloween kostymer njuter av en föreställning.
En liten flicka i blå rock gungar på en röd lekplatsleksak.
En man i kostym passerar en skivaffär.
En man går två pudlar på koppel i en stad.
Lilla flicka i blå klänning använder en rosa hula-hoop.
Ett lag hundar, och en kvinna som följer på en cykel.
En man spelar stålfat nära vattnet när folk passerar förbi.
En man i gul hatt har en färgglad uppblåsningshammare.
Tre personer går förbi en man som spelar flöjt på trottoaren.
Unga kvinnor bär en brun två stycke baddräkt bygga ett sandslott på en strand.
En familj ligger på verandan.
Tre personer tittar på marken nära ett bord och flera stolar.
Två små barn klättrar uppför trappan på ett plan.
Två hockeyspelare står och tävlar om pucken medan en målvakt hukar framför nätet.
Vandrarna klättrar upp för bergen.
En löpare får en vattenflaska från en kvinna i en töljacka som håller i ett paraply.
En dam och ett litet barn stirrar på sig själva i en spegel.
En asiatisk kvinna i en rosa tröja som håller rökelsepinnar.
Ett barn glider ansikte först nerför ett metallrör
En man håller i ett handtag i vattnet.
En grupp människor tittar på en liten bebis med blont hår.
En pojke i baddräkt som går i sanden mot vattnet
En man i lila skjorta, omgiven av människor.
En orange katt med svarta ränder på en strand.
Ungar som spelar basket i en gammal domstol.
En grupp människor går runt ett trångt område med smuts på marken.
Den bruna hunden fångar en boll i luften.
En grupp människor håller i sig när de rider på kollektivtrafiken.
Flera människor går nerför en flyg av stentrappor under dagen.
Tre pojkar leker runt en fontän på en kontorsbyggnadsgård.
Våt flicka i gul baddräkt ser över klippan till en simmare i vattnet.
En brun hund springer mot tre andra hundar.
En man stirrar på en annan man som observerar hans rakningsteknik.
En Toyota lastbil parkeras utanför en upptagen butik som renoveras.
Det finns en stor gul grävsko mitt på gatan.
En man i en vit tank övredel med hjälp av en bärbar dator som sitter bredvid en hög pelare med en staty ovanpå.
En liten brun hund leker med en luddig toffel.
Två flickor i matchande rosa och vita klänningar och två mindre pojkar i matchande svarta och vita skjortor.
En kaukasisk man i svart t-shirt håller upp två pinnar.
Ett barn i en boll grop och ett litet barn som leker nära fötterna på den person som tar bilden.
Tre män är tillsammans, två sitter och en står.
En kvinna med röd mantel ska klippa sig.
Damen i den svarta skjortan lagar den andra damens hår.
En kvinna klipper en annan kvinnas hår när hon ler mot kameran.
Damen bär en blå skjorta från brandkåren.
En man i en blå skjorta som bär glasögon använder en tunn pensel för att måla på en stor duk.
Folk går nerför en gata förbi en skivaffär.
Benen och mellansektionerna av två personer med skateboard.
Ett nyfiken barn ses njuta av en projektor.
En man i lila får sin frisyr med en jättestor torktumlare vänd mot honom.
En man som sitter och läser på tunnelbanestationen.
En fullt klädd ung kvinna kör en stolpe ner i en simbassäng.
En ung pojke visar upp sig medan han går sin vita hund i ett område.
En pojke håller fast vid och springer tillsammans med en karusell.
En blond dam med solglasögon ler.
En stor lägereld på natten med flera personer som sitter runt den.
Två arbetare i orange väst utför sitt jobb.
En grupp män är klädda i gamla militärdräkter och bär instrument som i en parad.
En man hänger från kanten av en sten medan två andra fångar honom.
Hunden simmar genom vattnet mot vattenfallet.
Den lyckliga bruden och brudgummen väntade på att fotografen skulle fotografera dem.
Svart och vit hund i vardagsrummet står på bakbenen.
En grupp tjejer sitter i dansstudion.
En flicka som bär en blå kort och gul skjorta uniform kastar en gul softball medan en flicka i en svart och röd kort uniform och röd hjälm körs.
En ung flicka svänger på en bakgård.
En grupp barn leker på gatan där vatten sprutas.
En flicka i röd skjorta gråter utanför.
Två hundar på koppel anstränger sig mot varandra medan deras ägare går ifrån varandra.
Den lille pojken har en fjäril på sina smutsiga händer.
En kvinna i grön tröja sitter ner med en tennisracket på väg att träffa en tennisboll.
Man bär huvudduk som griper tag i ett träd i djungeln.
Ett barn i randig skjorta leker glatt bland några vattenfontäner.
Män sitter i trappan när en kvinna går förbi.
Svart hund med röd krage klättrar över staketstolpar.
Ett barn klädd som en pirat ler.
Två hundar springer bredvid varandra på gräset.
En man får lufttid på sin Wakeboard.
Två hanar sitter på en docka, varav en spelar gitarr, och ytterligare två står framför dem.
Två barn spelar ett spel nära ett scenområde.
Kvinnan i blå jacka och kvinnan i denim outfit med en grupp på ett berg.
En äldre man, som bär vit hatt, sopar en parkeringsplats.
En Veterans Parade med tre flaggbärare som visar upp sina flaggor.
En man på en lastbil dekorerad med flaggor och bunt.
En maskerad man i halloweenmask tittar på en kvinna.
En kvinna i svart blus som spelar kortspel.
Två honor, den ena blå, den andra svart, leende och skratt
En tjej i jacka på en säng.
Många människor är på stranden, nära en byggnad med flaggor som flyger.
Svarta hundar hoppar i poolen till en hand.
En man som bär en grå militärskjorta med medaljer och en ljusblå mössa med guld på viftar med armen.
En person vid ett bord, klädd i svart kostym.
En äldre herre, som bär t-shirt och shorts, vänder hamburgare på en stor gasgrill i rostfritt stål.
En mycket glad sångare i en extravagant outfit.
En kvinna som bär en skyltdocka går nerför trottoaren och pratar på en mobiltelefon.
Ett barn står ensamt och håller i en röd ballong och tittar in i en mörk insida.
En man som kör nerför gatan i en gammaldags brandmotor vågor på åskådare under en parad.
En gammal man med mustasch sitter ner och håller i en pistol och ler.
En kvinna som bär en röd duk på huvudet passerar framför ett blått skjul medan hon går nerför gatan.
En kvinnlig hejaklacksledare i en glansig blå cheerleaders outfit hoppar över scenen medan han uppträder.
En kvinna bär djävulsdräkt och poserar framför en fontän.
En grupp av DHL anställda poserar på parkeringen för ett fotografi.
Tre personer går på en stig mitt på dagen.
En servitris som pratar med en man på ett café.
Ett barn, som bär ett stängt blått paraply, går med ett annat barn som är under ett gult paraply, på en lerig stig.
En clown ler för en bild under en parad.
Två personer höjer armarna på en snöig kulle i bergen.
En kille i svart skjorta som står bakom disken i en affär.
En man sitter på en laptop, medan två män (en sitter, en står upp) möter varandra i bakgrunden.
En hund med en sele och en leksak munnen.
En kinesisk man som bär en traditionell kinesisk rishatt bär en balanserad börda över axeln med hjälp av en lång käpp.
En kvinna målar en kopia av en bild hängande på väggen.
Fyra sportfantaster går tillsammans med soppåsar på huvudet som läser C U B S.
Två män i vita uniformer med svarta bälten tävlar i en kampsport turnering.
En grupp människor marscherar i en parad på en solig dag guidar en Oscar den Grouch float.
Man skär tårta på en rosa matta.
En katt sitter på ett piano bakom öppen arkmusik och en glaslampa som är på.
En man med en röd fluga som sjunger ett solo med en full herrkör i bakgrunden.
En militär man som spelar trummor från America's Corp Fort Lewis i Washington medan han är i en parad
Den mest fantastiska fritidsaktiviteter utomhus camping.
En liten flicka med blont hår och blå ögon bär en tröja medan hon sitter bredvid en varm eld.
En man som skär en tårtbit på en kontorsfest.
En man i brun rock bär hjälm och cyklar medan han bär två plastpåsar.
En man i röd kostym står nära andra.
En kvinna i röd hatt och klänning sitter ensam på en parkbänk.
En man skrattar medan han bär en vit skjorta.
Medelålders kvinna som bär en vit solhatt och vit jacka, lägger handen i en mans byxficka.
Någon sitter på en gul motorcykel.
En yngre pojke är hos tandläkaren som håller någons hand.
En man rör vid en tavla på en vägg.
En dam och en man som knäböjer och håller i ett snöre medan en annan kvinna tittar på dem.
En man i gul skjorta skär sin födelsedagstårta.
En man i svart rock och blå skjorta pratar på sin telefon inomhus.
Ungdomar sitter på klipporna bredvid sitt fritidsfordon.
En man med en tatuering som håller en mopp nära en spelbutik.
Två man, en i baseballuniform kastar en boll.
En stor grupp människor som tittar på eld fungerar tillsammans.
En person i uniform står och deras skugga kastas bredvid dem.
En liten flicka är på ett baseballfält där en äldre man ger sig av mot publiken.
En gammal man i vit hatt sover vid en fiskebrygga.
Besökare färdas längs en bergsväg när de går längs ett säkerhetsstängsel.
En god samarit drog ut en extremt berusad man från gatan på trottoaren för att undvika att han blev överkörd.
En kvinna tittar i ett teleskop för att titta på något riktigt litet, troligen något slags vetenskapslabb.
Fem personer, klädda i mörkblå skjortor, ger en presentation utomhus.
Ett barn på stranden begravde sig i sand med bara huvudet blottat.
En kvinna som pratar med en grupp om tre andra kvinnor.
En flicka med ansiktsfärg på, som bär en röd skjorta målar en bild.
En kvinna ser ut som en man som hindrar en ung pojke.
En kvinna med glasögon och en gul skjorta håller ut handen.
Två killar på en strand som håller en tredje kille i armarna och vristerna.
En grupp unga män begravs upp till bröstet i sand.
En kvinna och ett barn går på en lövfodrad trottoar, på väg mot två människor ridande hästar.
Människor går förbi byggandet som sker i en stad.
Två män med väskor springer åt samma håll.
En man som håller en walkie talkie framför en öppen grön låda med kontroller i den.
En ung man i slips, kör på sin cykel.
En blond-hårig man klädd i mörka färger sitter bredvid en kvinna klädd i grönt och bär en svart basker.
En grupp män städar upp skräp.
Den leende kvinnan i den röda hjälmen håller utomhus ett mycket långt rep.
Folkmassor som dansar under en gatufestival.
En man och två små barn spelar musik för en grupp åskådare.
Tre män i ett vardagsrum har en diskussion.
En man som kör en grön jeep går över stora stenar.
En kvinna med tung makeup står bredvid ett rött ljustecken.
En hund fångar en frisbee när den hoppar på gräset.
Crowd samlas för att lyssna på ett band
En man som går över en korsning med långt hår, en grön huva och en ryggsäck.
Blond kvinna som sitter i en vit klänning.
Kvinna i vit bikini topp och blå shorts med kropp av vatten i bakgrunden.
Många cyklister tävlar längs en grusväg.
Två små pojkar, från midjan upp, i en kampsport match, en levererar ett slag och den andra blockering.
Två barn med gula bälten duellerar i en kampsport klass.
En gravid kvinna sitter vid ett restaurangbord och smeker sin mage.
En man med röda byxor på väg mot marken.
En grupp små barn, pojkar och flickor, spelar fotboll.
En ung pojke klädd i blått och vitt sparkar en fotboll.
En grupp människor bildar en procession, flera av dem håller skyltar med fotografier på dem.
Pojken i röda badbyxor hoppar på sanden.
Två asiatiska barn sitter i stolar på gatan på sommardagen.
En man svingar på ett rep ovanför vattnet.
Det är en man som svänger av ett rep som svingar in i en sjö.
Publiken på en match i LA intar sina platser.
En grupp frivilliga som arbetar med barn för att göra en leksakskörning utanför en leksaker r oss för barn i nöd.
En kvinna i svart fotograferar.
En liten pojke i baddräkt går över ett avloppsnät medan vattnet stänker på honom.
En svettig, tatuerad man spelar gitarr.
En fågels syn på fyra personer som står mitt i höga klippor.
Människor står eller går nära järnvägsspår.
En man i lila skjorta som kör en röd cykel.
En man ger en pojke high-five utanför en frisersalong.
Fyra barn, två flickor och två pojkar på äventyr i en kanot.
Människor med skyddsvästar står i ett fält med spadar.
En man i gul väst röker och arbetar på ett fält.
En man i tunga vindjackor som går genom ett fält.
Tre män i skyddsvästar arbetar längs en väg.
Två män i blå uniformer och grön väst.
En man kör en bit jordbruksutrustning på ett fält.
Tjejer försöker träffa bollen under en volleybollmatch.
Två hundar springer genom vatten med ett rep och röda flyter i munnen.
Två män tittar ner från byggnadsställningar.
En man i svart keps och blå skjorta letar efter guld.
En man i grön skjorta som slätar ut våt betong.
En äldre asiatisk man står bredvid ett stort fat ris.
En kvinna sitter bredvid en hink samlade musslor.
En man i svart skjorta spelar slagverk på en uppsättning tomma fem gallon hinkar.
En kvinna som säljer blommor i gathörnet.
En lång man och en kortare man som går och pratar, bär samma sandaler.
Två män fyller i papper till en man i röd skjorta som ligger bakom disken.
Ett band uppträder på scenen medan publiken höjer händerna och klappar.
En man står under en stor klocka.
Två män står i mörka kläder på en busshållplats, en läser tidningen.
En blond kvinna i jeans läser på en bänk.
En liten flicka i rosa klänning som gråter.
Män njuter av en smörgås på en gatumässa.
En stor, svart hund med något i munnen kommer ut ur en vattenpöl.
En man och kvinna som bär Musse Pigg öron i en publik.
En ung man sms:ar medan han står framför en affisch.
Två unga män står på trottoaren och pratar med varandra.
En svart man med en blå skjorta och en bling som stirrar in i kameran.
Kvinnan står mot väggen fylld med gamla annonser med en kort vit skjorta med jeansjacka och kjol.
En svart hane lutar sig mot en vägg med en vattenflaska.
Två långhåriga små flickor sitter på en plattform.
En kvinna i blå kläder drar en katt från taket på en bil.
Många människor går genom en fullsatt utomhusmarknad.
Två arbetare i sina hattar och skyddsvästar står nära ett gult betongblock.
En manlig trummis och en kvinnlig sångare på en föreställning.
En man i svart kostym och halm hatt håller en tennisracket som om det var en gitarr.
En fattig kvinna i sjal gräver efter stenar.
En man är böjd med utsikt över något på en stenig strand.
En kvinna som ger en kopp till en afroamerikansk man.
En man i svart skjorta som säljer frukt på marknaden.
Indiska damer dansar framför publiken
En man i bakgrunden som ska rulla en död med armémän och en död i förgrunden
En ung kvinna utför en balansstrålerutin framför åskådare.
En grupp människor står framför ett tåg.
Crowd shuffles förbi öppning i gammal struktur.
Två män klädda i vita skjortor knappa ner skjortor, vita hattar, med blå halsdukar bundna runt halsen
En man står utanför på ett café.
Folk står framför vattenmeloner på sidan av gatan.
Tjejen sitter i eld för en show
Två unga flickor bär baddräkter och står under fallande vatten.
En svart och vit hund springer i några löv.
En pojke i en renässansmässa kostym står vid bilar parkerad på gräs.
En svart hund och en brun hund som slåss.
En kvinna löder en bit metall som en man tittar på.
En ung man klättrar uppför ett berg, en annan följer nedanför.
En pojke gör ett hjul på en klippa.
En äldre herre tittar ner på sin öl.
Kvinna i vitt i förgrunden och en man strax bakom promenader med en skylt mot John's Pizza och Gyro i bakgrunden.
Lite tåg rider med familjen.
En kvinna rör om i innehållet i en gryta.
En stadsgata städas av en man i ett grönt fordon.
En grå hund utforskar ett fallet träd i skogen.
Fyra kvinnor som delar en måltid skrattar tillsammans.
Mannen i grön skjorta och last khakis står bredvid en grön jeep.
Tre flickvänner sitter på en mörk teater.
En äldre man kör en kärra med en älskad mans minnesbild nerför gatan.
En kvinna i grön väst tar en bild av en häst.
En ung pojke med röd skjorta står på gatan med armarna öppna.
En man som håller fast en liten flicka på en cykel.
En man i svart skjorta och en liten flicka i orange klänning delar på en godbit.
En man, som sitter, serverar mat till en liten flicka.
Kvinna och äldre man går sida vid sida på löpband i ett fitnessrum.
En kille sjunger in i en mikrofon.
En kvinna skyddar sina ögon från solen när hon går på en gata.
Folk går runt på en fullsatt marknadsgata.
Ett par i jeans promenerar nerför en gata som ligger i anslutning till ett område som blockeras av med orange nät.
Två flickor ligger i sängen med två små hundar.
En man och en kvinna poserar för ett foto bredvid ett klädställ.
En klättrare skalar en bergsklippa.
Två kvinnor som bär vad som verkar vara flygvärdinna kläder och solglasögon viftande inuti en byggnad.
En man står framför en prins St. Cafe.
Liten flicka i röd, vit och svart klänning ser på stora silver klot.
De små barnen klappar en gris
En hund går på en röd planka med ett blått räcke.
En äldre kvinna i en Burberry-rock, äter.
En kvinna i svart med en solbränd kostymjacka står på ett podium och talar till en publik.
En ung flicka som springer nerför en gata.
En man i slips spelar gitarr medan en välklädd kvinna tittar över noter, möjligen för att sjunga.
När jag har utsikt över staden hämtar jag min gitarr på grund av inspirationen.
Ett blond barn springer nerför ett fält och tungan sticker ut.
En kille läser en bok när han sitter framför ett piano.
En person raderar en båt över en stor vattensamling.
En hund på en strand som släpar ett föremål
En mor vaggar sin skolelev i famnen.
En kvinna sätter upp en stege för att måla taket.
En person på en cykel har en vit hund i koppel.
En kvinna med glasögon ger en presentation till två kvinnor som sitter ner.
En kvinna får hjälp av kvinnan bakom disken.
En man i grön skjorta håller fram en urtavla för en kvinna i rosas uppmärksamhet.
En manlig vakt står bakom en annan man i en mönstrad tröja.
Två killar, i svarta skjortor, som röker utomhus.
En kvinna i svart bläddrar genom sidor i en bok i ett bibliotek som en flicka i vitt med hörlurar ler.
En kvinna som hjälper en annan kvinna med en hemsida på en dator.
Två barn faller huvudet först i en färgstark boll grop medan ett tredje barn klockor.
En detaljhandeln professionell pauser samtidigt interagera med kunder.
Tre hundar springer runt i gräset med skog i bakgrunden
Barn och vuxna leker i grunt vatten i en stad.
Groom bär svart och grå smoking och brud bär en vit klänning är beströdda med blommor.
En lycklig, vacker brud som kliver ur en lyxbil.
Man cyklar genom diry cykelbana bär vit hjälm och handskar
En grupp människor som har samtal på en restaurang.
En Houston basebollspelare har fångat en boll och kastar nu bollen mot en annan lagmedlem.
Tre personer på scenen sjunger och spelar instrument.
Tre personer handlar i en ö i en utländsk livsmedelsbutik.
Fyra pojkar hoppar in i en inomhuspool.
En liten vit hund klättrar över en stock.
En dam som sätter upp flerfärgade bollar i en tramption.
Två män, båda bär ljusgula västar och jeans, arbetar på ett tak.
En man i vit utstyrsel spelar ett elektriskt tangentbord.
En man i en floppig hatt och ljusa gula shorts står i lera.
En man talar in i en mikrofon.
En äldre man går nerför trottoaren med svarta shorts och en vit skjorta.
En rödhårig kvinna som pratar i telefon medan hon klappar en brun och solbränd hund.
En man står under en valv nära Wendys restaurang.
Ett gossebarn som håller en boll stående på trottoaren.
En väg är blockerad och polisen är på väg runt den.
En grupp ungdomar sitter och pratar.
En vanlig kille som tar en drink i en asiatisk bar.
En hund skakar vatten av sig själv.
Två hundar drar på en rosa och orange boll från motsatta ändar.
En man i tillfälliga kläder håller en presentation.
Ett nyfött barn sover på sin sida efter en lång dag.
Två herrar är mitt i en datorklass.
En kvinna som bär en T-shirt, shorts och sandaler, är minigolf framför blommor och en gångväg.
Fyra män går på gatan i kallt väder
En flicka står på gatan, och den andra hukar sig och tittar på något på marken.
Två personer sitter framför datorer och ett stort mörkt fönster.
Folk rider och rodder en båt nära kusten.
Två män, en med en svart sopsäck.
En man i tröja lägger en sopsäck över en brevlåda.
En man i svart skjorta och baseballmössa som plockar upp skräp på en tom tomt.
Ett barn leker med mat medan det sitter i en barnstol.
En man sitter på en röd duk på marken nära en blå stolpe.
En grupp tonårspojkar som går längs vägkanten med en sopsäck.
En flicka och en pojke sitter bredvid varandra i ett fordon.
En man med visir och blå topp har kastat en frisbee i fjärran.
En kille som ska kasta en frisbee.
En man kastar en blå frisbee mot ett frisbee golf mål.
Två män packar munkar i plastfolie.
En pojke i en grå tröja kastar en påse skräp i en grön container.
Män och kvinnor som äter som en kvinna arbetar på en dator.
Två asiatiska kvinnor håller upp en delvis fylld sopsäck, ler.
En svart man som bär sönderslitet tyg.
En ung man tar en påse skräp till sopcontainern, efter att ha plockat upp skräp på gatan.
Ett par går på en trottoar längs en strippklubb.
En man som bär en grön tanktopp och en vit hatt som sjunger in i en mikrofon.
En ung man i en färgstark kostym sjunger in i en mikrofon.
En man kastar en sopgubbe i en container medan en annan håller locket.
Män i färgglada skjortor visar kamratskap efter en cykeltävling.
En pojke flyter med hjälp av en brun apparat i en vattenförekomst.
En grupp människor i hårda hattar bygger ett hus.
En grupp byggnadsarbetare som bygger ett hus.
Tre män bygger ett tak.
Fyra barn läser ett recept i ett professionellt kök medan ingredienserna läggs ut på bordet.
Två personer med cyklar stående framför en byggnad.
Det finns en grupp barn som får sin bild tagen med presenter.
En fiskare har sin fot fångad i sitt nät.
En skjortlös man med ljusblå shorts och en keps står framför en båt.
En man står i vattnet och tänker på något.
Två män klädde upp sig inför en stor tillställning.
En man sjunger och spelar en vit gitarr.
En man som går medan han håller ett litet barns hand.
En tonårspojke utför ett stunt på sin skateboard i en skatepark.
En äldre man står bredvid en uppvisning av träbrickor.
Coeds sitter på ett picknickbord i sten och äter lunch på gården.
En man står nära en gata i kostym med en skylt som säger "Sluta våldta min fru!"
Folk åker skridskor på en rullskridskobana.
En pojke med rött hår håller upp en glasstrut för en äldre man att provsmaka.
En ung pojke leker i en bäck säng
Människor i ett mörkt rum som har väggar upplysta av grönt ljus och en person håller upp sin mobiltelefon.
En man med skjorta och slips på toppen av ett hissschakt.
En man som pluggar in en tråd medan han håller i en gitarr.
Två män använder verktyg som skär in i en grön trailer.
En far och hans son skär en tårta under en middagsbjudning som hålls på deras residens i Texas.
Två män står och en har en slang.
Våt svart och vit hund med svart näsa skakar av vatten.
En blondhårig kvinna går en hund nerför gatan i flip-flops.
En man i blå skjorta går och håller en ung pojkes hand utanför i en trädgård.
En pojke står i vattnet nära en frisbee.
En kvinna sitter med fötterna i en grund pool och tittar på en valp.
En man med en blå mask som läser en bok.
En svart och vit hund som bär en sele slickar en brunett i glasögon.
Kvinna i grön topp och blå jeans bowling.
En man med en cigarett i munnen kör motorcykel.
En grupp barn i blå kläder står vid en grind.
Två män i vita skjortor som jobbar i en gammal byggnad.
En gatuscen med mötande trafik, inklusive bilar och motorcyklar.
Två kvinnor bär grå t-shirts, en håller två bruna papperspåsar, lämnar en kartlagd buss.
En kvinna i en tank-top, skära en annan kvinnas kläder.
Ett barn med brunt lockigt hår som njuter av en drink.
Stor utrustning som rör sig på marken i arbete.
En man i hård hatt sköter en grävling.
En brun hund i en kanot tittar ut över stilla vatten.
Tre män i vitt målar räcket på piren blått.
En grupp människor som sitter på ett däck.
Folk har ett samtal och en vattenflaska föll ner på marken.
En pojke i blå och gröna byxor ligger mot en vägg.
En brun hund står framför några växter.
En man brottas med en tjur medan åskådare tittar.
En äldre kvinna som köper schampo och balsam i en butik.
En fotograf fotograferar blommor.
En bergsklättrare lutar sig ut från en klippa mot en djup blå himmel.
En man och en kvinna i glasögon blåser bubblor.
En grupp unga män brottas och horsar runt i en smutsig grop.
Kvinnorna håller en bild av ett barn som ligger på marken.
En man i vit rock skär kött med en mycket vass cleaver.
Det ser ut som körträning i en äldre utsmyckad kyrka.
En man går nerför gatan en höstdag och sparkar löv i luften.
Mannen i orange skjorta håller tal.
Två barn leker med en fotboll på gräs.
En liten rödhårig pojke spelar Whack Em!
En hund hålls i koppel av en kvinna i vita skor.
En man som rakar sig med rakkniv.
En kvinna äter en sallad i läktaren på ett arenaevenemang.
Folk letar efter sina platser på en stadion.
Två småbarn äter majshundar i en liten vagn eller soptunna.
Cyklister, en kvinna som knuffar ett barn i en barnvagn, och människor som sitter i en park.
En ung pojke i blå skjorta står bredvid en kvinna som sitter på marken.
En kvinna sträcker sig in i en låda med godis medan en man står i närheten.
Flera människor ser ett kvinnligt rockband uppträda på en scen full av gula banderoller.
En kvinna lyssnar på bandet på scenen.
En äldre kvinna som ler, i en blå rock, med sin hund.
En man duschar i ett hem utomhus duschanläggning.
En man i blå skjorta tittar upp på ett barn med röd randig skjorta och blå jeans.
En man i en kvinna i ett hus umgås glatt.
En man städar sin trädgård med en lövblåsare.
En man och en kvinna tittar uppåt på ett kvarter.
En långhårig man spelar bandspelaren och en mås sitter i närheten på en vägg.
Två personer springer på stranden av en strand
En liten pojke som ser barn som bror får en hennatatuering.
En man i grå skjorta gäspar.
En kock som arbetar på en spishäll som är täckt med krukor och olika redskap.
En pojke gömmer en fisk medan en flicka pekar på fisken.
En frisör i svart skjorta skär försiktigt en ung pojkes hår.
Två snorklare befinner sig i ett mycket blått hav och simmar med en orange boj.
En kvinna i förkläde och vit skjorta står bakom ett fullt buffébord, medan en man är böjd bakom henne.
En grupp äter lunch på rasten.
Två män sparkar i en ring, en man slår den andra.
Folk står i en rörig gränd.
Två små asiatiska pojkar poserar för kamera i ett grönt inhägnat rum.
En grupp människor sitter i en cirkel och roar sig.
En liten gammal kvinna klättrar ut bakom den blå dörren och tre par sandaler i plast.
3 personer i en liten stuga eller hus.
Ett litet barn hålls ovanför en mans huvud när hennes hår flyger i luften.
Två män som cyklar på motorvägen.
Det finns grupper av flickor från olika etnicitet gör barn hejarklacksrörelser i ett gym på en matta.
En man i khakibyxor står på en soptunna och kramar om en stolpe.
En grupp människor hoppar ner i en sjö unisont.
En hund som dricker ur en vattenspik.
Ett barn knuffas av en stor våg medan han håller i sin gula surfbräda.
En utexaminerad student i kläder talar med en professor.
En vit flicka svingar ett svärd.
En obekväm tjej som tittar ut genom ett fönster på gatan utanför.
Två män vandrar med ett litet barn nära några intressanta form klippformationer.
En medelålders man som bär röd hatt fiskar.
Två pojkar står på sanden bredvid en vältad stol.
Pojke med blå handduk och vit hatt som håller goggles och en snokel.
En pojke som simmar och bär glasögon.
Ett barn som tar en paus från att leka och äta glass.
Någon tar av en Green Bay Packers-fotbollsspelare.
En kvinna med en budbärare väska cyklar.
En brindle-belagd hund morrar på en hoppande brun hund med lila krage inuti en park inhägnad.
Tunga maskiner i bruk på en fabrik.
Två pojkar är fast i ett träd och svänger över en tråd.
Fyra kvinnor arbetar tillsammans för att laga mat.
En asiatisk man ligger på ett kaklat golv med två barn och använder gamla kläder till kuddar.
Tröjlös man balanserar på ofärdigt tak.
Två män i skottsäkra västar vakar över en folkmassa vid några vita tält.
En liten pojke som spelar fotboll i parken.
En liten pojke i en blå skjorta som sparkar runt en fotbollsboll.
En man som går in i skuggorna.
En grupp soldater hukar sig över en eldgrop med köttkokning på grillen.
Äldste man arbetar med ett projekt i sitt hem verkstad.
En ung man röker en cigarett medan han håller i en maroongitarr.
En äldre man är utanför och bär på växter.
Två barn i badrummet, en står medan den andra läser en bok och använder toaletten.
Två asiatiska män i mörka kostymer som pratar.
En man klädd i svart och vitt använder ett vasst verktyg för att hugga trä.
Två personer på en båt tittar på solnedgången.
En flicka klädd i blå och bruna väskor stående i slutet av en tunnel.
Tre fönsterbrickor i blå uniformer fungerar på byggnadsställningar.
Två unga män leker utanför nära en gyllene staty av Ghandi.
Två hundar leker med en leksak utomhus.
Två män tävlar runt ett grusspår på cyklar medan en handfull åskådare tittar bakom ett staket.
En kvinna som sitter i en park och pratar på en mobiltelefon.
Tre personer står nära tre flerfärgade varmluftsballonger.
Sex mycket färgglada varmluftsballonger gör sig redo att flyga.
Pojken håller en basketboll på en basketplan i trä.
En pojke dribblar en basketboll i gymnastiksalen.
En ung pojke i rörelse framför krukväxter och en beige vägg.
En ung kvinna med en blå hjälm som klättrar upp för en sten.
En man som bär vit t-shirt och shorts är att klättra med andra människor som bär blå hårda hattar.
En dam blåser upp en otrolig hulkleksak.
En person i en fallskärm med en amerikansk flagga fäst vid honom.
Någon är fallskärmshoppad och nästan rör vid marken.
En ung flicka i randig skjorta har en elektronisk ljudmakare som hon byggde själv.
En man fallskärmshoppar bredvid ett jetplan.
En erfaren fotograf knäpper fotot trots att han är nertyngd av all sin utrustning.
Små barn har kul när de spelar säckhoppning i parken.
En grupp barn har kul i säcklopp.
Baby sover i sin bilstol.
En man i grå jacka och vit skjorta lutar sig mot ett räcke och pratar med en annan man.
En medelålders man som kör sin svarta motorcykel genom ett kvarter.
En man i svart skjorta åker förbi en bänk i stan.
Två män filéer en fisk i ett handfat medan andra tittar.
Folk sitter på trappan längs vattnet och fiskar.
En kvinna som hänger på en flotte.
En kvinna med kort blont hår reser sig från en stol som en annan kvinna i en bourgogneskjorta skrattar.
En kvinna som bär en rosa skjorta använder träningsutrustning.
Tre personer går på en regnig natt på en gata i Kina.
En man som bär shorts och ingen tröja hukar sig.
En cykel står parkerad framför en butik som har en stor orange skylt.
Förbereder en fiskmiddag för familjen.
En pojke med blå hatt pekar mot en skål full av kork.
En kvinna håller i ett barn medan ett annat barn står vid hennes sida.
En pappa och hans pojkar är ute som en familj och sköter familjesysslorna med sin boskap.
En man med hatt lagar grill.
Tre kvinnor i olika åldrar i vita klänningar sitter i en dammig glänta framför träd.
Passagerare som åker järnväg genom stan.
Två kvinnor i uniform står på sidan av vägen när en kvinna i vita cowboystövlar går förbi.
Jag tror att byggnadsarbetet pågår här.
Fem vandrare färdas en torr, skrubbig slätt mot snöiga toppar i bakgrunden.
En grupp barn håller ballongdjur.
En flicka i grön jacka knäböjer och tar en bild av en annan flicka som står upp.
Man i vit polo t-shirt med glasögon spelar en röd gitarr.
En skjortlös man som dyker ner i en inhägnad grön pool medan det finns en skog bakom honom.
En kör som sjunger för församlingen i kyrkan.
En man sitter på en bänk framför några lila växter.
Två personer med cykelhjälmar chattar på en bänk.
En man i orange rock stod på en stege och inspekterade en enorm metallbehållare.
En påträngande kvinna klättrar över ett stängsel.
Medborgare njuter av en snöig dag med påminnelse om sommaren i bakgrunden.
En tjej i overall gör en snöängel.
En man sätter rakkräm på skägget medan han tittar i en spegel när en annan man står i bakgrunden.
En man iakttar antikviteter i en affär.
Två kladdiga gula hundar som leker på ett tufft sätt.
Flera byggnadsarbetare som bygger en parkeringsplats.
En grupp pojkar spelar flaggfotboll medan några åskådare tittar på.
Det finns många människor på gatan.
En skara män i uniformer bestående av blå toppar och vita byxor går.
Mannen installerar kakel på badrumsväggen.
Två killar installerar kakel i vilket är kanske ett badrum
Folk trängs in på en gata i en asiatisk stad.
En grupp människor står på sidan av vägen med en orange buss bredvid dem.
Fyra asiatiska människor paddlar kanot i tre kanoter.
En grupp turister ombord på en liten och färgstark båt i vattnen i ett sydostasitiskt land.
En folkmassa samlades runt en man som bar en röd japansk mask.
En person med ett randigt rör som står mitt i en folkmassa.
En leende person med jacka och stövlar hoppar i en stor pöl.
Tre personer vandrar uppför ett berg med en flod och andra berg i bakgrunden.
En kille och en pojke rider på en skateboard tillsammans.
Två dachshunds springer i gräset med en blå boll.
En apotekare är på jobbet och fyller på recept.
En flicka sjunger i en mikrofon medan andra tittar på henne.
En brun hund som leker med en tennisboll
Fyra killar i en bil med en i mittsätet vände sig bakåt och tittade på kameran.
En man håller upp en plastburk inomhus.
Tjej i röd rock, blå huvudduk och jeans gör en snöängel.
En grupp flickor som har en studiefest.
Person i huva tröja som skymmer ansiktet sitter bredvid en nyskuren stock.
Män som har en trädsnideritävling.
Två män i neongula skjortor sågade ivrigt en stock på mitten.
En grupp tonåringar pratar nära en cementvägg.
Kvinnan står framför en stendamm och bär en röd skjorta.
En man i gult hi-viz griper tag i en träbräda.
Två män sitter på en järnvägsslips och visar kameran något i handen.
En man gör kringlor i köket.
En grupp barn står på scen inför en publik redo att uppträda.
En kille knuffar en vagn full med vatten i väskor på resenären.
En kvinna i lila klänning inspekterar ett stort tygstycke.
En kvinna sover medan hon sitter på en parkbänk.
En man i en hård hatt står ovanpå en hög med spillror.
En orientalisk kvinna på en fullsatt gata som pekar.
En brud och någon från hennes bröllopsfest, klädd i en mörkare klänning, går på stranden.
En silverstaty av män på cyklar.
En kvinna derssed i en svart tröja, handskar, hatt och en halsduk sitter på stranden nära ett stenblock.
En liten pojke står på en kamrat bredvid en båt.
En gymnast i en blå leotard gör ett handstöd på träningsgolvet.
Ett barn i gröna skor som stirrar ner i ett avlopp.
En vit man i gul skjorta som säger "Glass Collector" drar mycket hårt på ett mycket stort rep.
En pojke i kamouflagebyxor och en orange skjorta har hatten baklänges.
Många människor på gatan framför stora byggnader.
En brun hund springer genom grunt vatten med en käpp i munnen.
En man i randig skjorta ser en tunnelbanebil köra förbi.
Vissa män lagar nåt mitt på gatan.
En skallig man med färgade tatueringar på armarna stannar i skogen med två hundar.
En man står på toppen av en sten medan han tittar på en cykel.
Ett barn i orange leker med en snöboll utanför.
En person går uppför en snöig kulle
En man i shorts står på en klippa och tittar ut över utsikten från kullen.
Den bruna hunden går genom blommorna.
Kvinna som bär blå bikini nedredelen och blå sportbehå kör på en atletisk bana.
En kvinna och två män i ett klassrum.
En brunetttjej med glasögon och en blond tjej pratar ute på ett fält.
En brun hund hoppar upp för att fånga en tennisboll.
Fyra män (2 observerar) med hjälmar gräver i marken.
En gammal kvinna väver ett tyg.
Vilken vacker dag för en ensam snorklingsexpedition.
En brun hund och en liten tjejkyss.
En avlägsen figur går mellan träd med en lätt dammning av snö på dem.
En hund springer för att fånga en frisbee på AstroTurf.
En pojke i röd baseball utrustning gör en pitch, framför en trailer park.
En stor skara människor samlas på gatan.
Person som sitter i en stol och säljer varor utanför en byggnad.
Ett barn leker med en vatten pip utomhus medan resten av sin familj tittar.
En kvinna med kort blont hår håller sin violin och båge.
En man går nerför ett snöigt berg.
Två pudlar är i snön och en hoppar högt
Chefer på balkong tar en paus från arbetet
En stor grupp människor i en röd flotte bär röda flytvästar på floden
En man med upplyfta armar på toppen av ett berg.
Ett barn spelar en röd leksak gitarr och sjunger i flerfärgad plast mikrofon.
En man som paddlar i vatten.
Två män är ivriga att njuta av en läcker kalkon i ett stökigt kök.
En man förbereder en måltid på en köksdisk med tre skålar.
En skallig man med glasögon skär i en kalkon på middagsbordet.
En man med svart hår stirrar åt höger.
De lila fallskärmarna flyter från klippan mot det grå havet nedanför.
Fallskärmshopparen står på ett fält nära sin fallskärm.
En man sätter en kalkon på en grill.
En grupp arbetare bygger något.
Tre kvinnor samtalar under ett paraply, med en annan kvinna som sitter ensam på en bänk.
En man i blått som gör kung fu.
Fallskärmshopparen har en fågel som flyger med honom.
Två fågelhundar tävlar om att döda.
En man föreläser om en grupp människor i ett medelstort rum.
Ett barn som knuffar sitt yngre syskon i en barnvagn.
En tjej i blomklänning springer på sand.
En liten vit bebis sitter i en resväska.
En skara människor går, de är mestadels klädda i vitt.
En bild på två flickor som använder garn på natten.
En svart valp med svart krage sitter på gräset och lämnar.
En liten asiatisk pojke kryper fram på asfalt.
Ett barn som bär en mörkgrön rock som bär en leksak i en leksaksaffär.
Ett barn har en spelkontroll ovanför huvudet och skrattar.
En äldre man lägger en trälåda ovanpå en hög med trälådor.
En man som lutar sig mot skrivbordet och lyssnar på någon i telefon.
Det ligger en man på marken med en röd och vit hatt på huvudet.
Tre pojkar i ett trä-panelat rum, en inspekterar en båge.
Det finns tre män, som verkar vara identiska, som sitter vid ett skrivbord med den på slutet dricker från en kaffekopp.
En man pratar med en pojke i ett ledigt område.
En grupp unga vuxna kvinnor sitter i golvet och stickar.
En man knuffar en pojke på en lina.
En brun och svart hund springer längs en gräsbevuxen stig med en röd jacka.
2 vandrare är i vattnet försöker korsa.
En asiatisk man leker med sitt barn i en modern lägenhet.
En ung familj sitter på trappan och njuter av dagen
Vuxna och barn står och leker framför trappan nära ett skogsområde.
Två barn som står mellan två röda bilar.
En man sitter med en kopp kaffe och läser en tidning.
En man i vit skjorta som håller i en snöskyffel.
En brun hund och en svart hund är tillsammans i högt gräs.
Folk går i en stor pöl.
En man jobbar på bältros på ett tak.
Tre barn brottas på en blommig matta.
En man flyger genom luften när en ung flicka står på en soffa och slår honom i magen.
En arbetare som hänger i en hög metallstänger.
Här är en bild av en man som arbetar med ett byggnadsarbete.
Tre hundar springer över banan.
En dam i rött står mitt på gatan mellan linbanespåren.
En liten pojke dansar på betongen omgiven av vuxna.
Ett litet barn leker med en leksak framför en vägg.
En man och en kvinna är i stan och ler.
Solen skiner över snön och träden.
En läkare konsulterar en patient.
En stor publik och kamerabesättning möter en idrottsplats.
Det finns ett stort skelett bakom ett stängsel.
Ryttarna och hästarna tar en paus och vilar på fjällstigen.
Två små barn går nerför en trädkantad stig.
En grupp muslimska män ställde upp i bön i ett stadsområde.
En man håller och matar sina två små barn.
En man som bär en svart skjorta dammsuger gräset.
En liten pojke som drar en grön vagn i tröja och stövlar.
En manlig läkare mäter en kvinnas blodtryck.
Två hundar slåss på sand.
En liten flicka i en blå och rosa leotard går längs en bjälke medan en persons hand sträcks ut för att stödja henne.
En dam och en kille sätter sig ner och slår in presenter.
En barfota ung pojke tittar på kameran medan han svänger i en park.
Två bergsbestigare ler på bergssidan.
En man med ett mörkgrönt förkläde som står med händerna på midjan med en grill i bakgrunden.
Ett litet badkar sitter framför statyn.
En blond kvinna dansar en solig dag.
En man ger en annan man mat från en utomhusförsäljare.
Två gamla män använder Jackhammers på trottoaren medan folk går förbi.
Två barn, båda i röda jackor, leker på trappan utanför.
En ung flicka hoppar från en soffa och högt upp i luften.
En person i vinterutrustning är att cykla nära en korsning.
En hona med svart halsduk och hjälm som cyklar.
En person tittar ut genom fönstret på A-bussen.
En vit hund med falska horn på huvudet och en brun hund leker tillsammans utomhus.
En liten flicka klädd i rosa spelar hopscotch.
En kvinna klädd i svart klädsel och orange halsduk stående mot väggen bredvid kartan.
En grupp människor samlas vid ett träd.
På övervåningen, på ett café, äter en man och vid ett separat bord talar en annan på en mobiltelefon, medan en man där nere sitter bland kartonger.
En blondhårig pojke och en brunhårig flicka skrattar tillsammans medan de äter.
En kvinna i en ljus klänning som skrattar.
Två män lagar mat medan de står i köket
En person gör en vända mitt i fältet medan deras vän tar en bild.
Några unga män spelar basket.
Tre tävlingshundar springer ut från startgrinden på ett spår.
En brun hund som springer på en gård.
En asiatisk man i svart rock håller upp en liten fläkt av en buske med rök som kommer ut ur den.
En man skateboards nerför ett brant räcke bredvid några steg.
En mörkhyad man cyklar på en gata full av trafik.
En man ser på när en annan man stuntar på sin cykel.
En grupp vandrare som tar en kort paus.
En hund hoppar in i en simbassäng efter en anka.
Kvinnan bär rosa hatt och cyklar i parken.
En kvinna jonglerar sitt barn, handväska, pengar och mat från en marknad.
En flicka som är omgiven av andra människor tar en bild på en konsert.
En man i brun rock pratar med publiken.
En grupp motorcyklister sitter på sina cyklar på en gata.
En vacker dam sminkar sig i spegeln.
En man klädd i en klänning som går fram till en duk, åskådare tittar på
En svart valp som tuggar på en brun hunds hals
En äldre kvinna presenterar en tårta för en grupp barn.
En liten flicka går mot trappan där det finns en duva.
En brun hund jagar en vit hund genom det lummiga gräset
En gammal man, med grått skägg, rider sin cykel
Två små pojkar med brunt hår och en med blont hår.
Två poliser står i ett livligt gathörn.
En person på en strand i en grön hängglidare.
En kvinna klädd i svart och guld som tittar åt hennes sida.
En kvinna som ser fram emot att titta åt höger.
Två kvinnor i kjol går längs gatan.
En vandrare skuggas av tiden på dagen nära en öppen och trädfodrad vattenförekomst.
En man som står vid en röd bil och ett litet barn tittar ut genom fönstret.
En man som kastar ut en fiskelina i en bäck
En person går bland stor, vit geometrisk formad arkitektur.
En man vandrar på en bergstopp en molnig dag.
En kanot på väg mot en annan på en dimmig flodbank.
En man äter något och går nerför en trottoar förbi en stor röd och gul skylt.
En tjej som sitter på marken pratar på en mobiltelefon.
En östasiatisk kvinna sitter i vad som verkar vara en tunnelbanebil när två affärsmän står framför henne.
En kvinna har grönsaker utlagda på en display.
En målare hängande på sidan av en byggnadsmålning, med två hinkar fastspända vid sidorna.
En man i vit skjorta tittar på en gatuförsäljare.
Två damer som går på trottoaren och pratar med varandra.
Kvinnor som fjäskar över sitt nyfödda barn och sitt lilla barn.
En man och en kvinna som bär påsar går nerför trottoaren.
En pojke sitter i biblioteket och läser en bok.
En brun och vit hund håller en tennisboll i munnen.
En grupp människor i skyddsutrustning.
En kvinna med långt rött hår står i sitt vita kök och håller en svamp och ler till personen som tar fotografiet.
En grupp människor sitter på bryggan och dricker några öl.
Det finns tre män som har ett samtal på en social plats.
En hund springer i skogen.
Två kvinnor kramas i ett trångt rum där folk dricker.
En grupp människor i en byggnad.
En brun hund med hyreskontrakt springer med en person bakom hunden.
Två män som har ett samtal i en utomhus allmän plats.
En man med glasögon satte sig precis ner och är redo att äta sin hamburgare.
En ung man i blå skjorta äter en korv.
Två barn i rockar poserar med en snögubbe.
Fyra personer tittar genom ett stängsel på något.
Två leende unga män ligger i en grön papasan stol med en solbränna tröstar över dem.
En stor grupp människor samlas utanför.
En flicka satt vid ett bord och försökte göra ett pepparkakshus.
En man som tittar ut genom ett tågfönster.
Tre barn hoppar in i en pool med en palm i mitten.
Två barn i identiska kläder hänger på ett kedjelänkstängsel.
En pojke i pyjamas byxor hoppar på en röd soffa.
En man lagar korv klädd i typiska kockkläder.
En svart hund leker med lite is vid den frusna floden.
Folk går nerför gatan på en mässa.
En äldre kvinna cyklar i staden när en gul taxi är på väg att passera.
En kvinna som stod i en dörröppning och rökte en cigarett.
Mannen bär en halsduk, jacka och en pälsig hatt en snöig dag.
En pojke leker cricket.
En mamma är väldigt glad över att få hålla sitt nya barn.
En svart och vit hund hoppar i gräset.
Den svarta och vita hunden tillsammans med den bruna hunden galopperar utanför
En kvinna med hjälm som cyklar.
Två pojkar som spelar cricket, en kastar en orange boll.
Ett porträtt av en flicka och ett litet barn.
En man ser ner när ett barn sover i hans armar.
En flicka håller i en boll och pekar på en frisbee.
Skolbarnen bar uniformer av vita skjortor och marinblå byxor eller kjolar och gula namnskyltar.
Sju personer sitter vid bordet i metall fällbara stolar diskutera ämne.
Ett litet svart barn står på kanten av en vattenförekomst nära hinkar.
Ett medelstort barn hoppar från en dammig bank över en bäck.
Folk beter sig som om de väntar på svar från någon eller något.
En kvinna som bär en röd kjol går bredvid en stenmur.
En röd hund hukar sig i snön.
Ett litet barn dansar på en halmyta.
En pojke drar ett vilt ansikte medan han viftar med kokredskap i händerna.
Två tjejer som håller i drinkar och tittar på något på en mobiltelefon.
Ett litet barn i stickad mössa och rock har en snöskyffel i en snödriva.
En grupp människor tittar in i sina kameror
En man på en kajak kommer nerför ett rasande vattenfall
En man i en gul båt paddlar nerför grovvatten.
En liten flicka i lila klänning tittar ner på kameran.
En man ler i sin blå och gröna kajak.
Kvinna och en man som står tvärs över gatan från varandra på en korsning.
En man och en kvinna dricker på en bar.
En man på en parkeringsplats bredvid en röd lastbil lägger en låda i den.
Den bakre änden av ett djur vars främre ände är under jord.
En mustad man i vit skjorta befinner sig vid en monter som visar cigaretter och glasflaskor med olika läskedrycker.
Verkar vara en stor samling av människor som rappade i bourgognekläder.
Två män klädda med päls runt sig med hela näsor och hattar och solglasögon på.
Folk poserar för en bild i snön
En ung vit man, klädd i mörka byxor och en ljusfärgad t-shirt som spelar ett franskt horn i ett band.
En äldre man i en Hawaiisk skjorta som bär en stor bunt på axlarna.
Ett skadat fordon bärs av en reparationsbil på en nattlig scen.
Två små flickor ligger på gräset och ler.
Två män, utan skjortor på, spelar bordtennis
En man som bär solglasögon spelar gitarr.
En man med en svart skidmössa och ett rött och vitt pannband tittar i fjärran.
En barfota liten pojke sopar ett tegelgolv.
En hund med en tidning i munnen springer nerför en asfalterad stig.
Tre kvinnor sitter på en bänk och väntar på bussen.
En man i svart kostym surfar i havet.
Tre svarta hundar simmar i smutsigt vatten
En ung flicka som håller en tårta med ljus klädda i en tung kappa.
En brun hund går i vattnet.
En man i brunt och rött spelar golf inomhus.
En man vandrar på en grusväg högt över en stad.
En ensam vandrare på en grusvandringsstig med hatt och solglasögon på med träd i bakgrunden
Hiker står på toppen av en sten med utsikt över en stad.
Två män står nära en stor maskin.
Två män, klänningar i jackor och handskar, blåser löv.
Två män i arbetskläder står bredvid en artonhjuling utanför en stor fabrik.
Kvinnan och barnen står bredvid en staty av en ko.
En man i grön hatt tar ett självporträtt.
Tre vuxna med kall väderutrustning.
En pojke som bär svart går nerför gatan med händerna i nävarna.
Två flickor spelar på en skateboard på en gårdsplan.
En kvinna i röd rock och brun hatt och en man i svart skinnrock går förbi en gatuförsäljare.
Brunhårig hane som slappnar av i en ek.
Stor fluffig grå hund står i gräs framför en brun hund.
Mannen i gul usa-skjorta sitter utanför entrén.
Denna jordbrukare skär i sin skördade frukt med en machete att sälja på marknaden.
Fyra kvinnor på en bar som skrattar.
En grupp män och kvinnor som sitter på bås och dricker ut flaskor och glas.
En svart hund går över sanden.
Folk sitter vid långa matbord i ett tält vid något formellt evenemang.
En ung kvinna ser glad ut i vinterkläder medan det snöar.
En man och ett barn går längs stranden när en boll flyter i vattnet.
Ett orkesterband övar i en kyrka.
En liten pojke med grön skjorta springer på en klippavsats.
Två unga män säljer varor på en marknad.
Två tjejer hoppar på en studsmatta, en upprätt och den andra landar på ryggen, på en bakgård.
Folk står utanför och ser motorcyklar köra på en väg.
En äldre man i vit skjorta som kör motorcykel.
En person går förbi något blågrönt vatten medan han håller i en rail.
En grupp motorcyklister kör runt en parkeringsplats.
En man som ristar en pumpa i sina boxare.
En ung flicka som står bakom en Davidsstjärna.
En person ligger halva under en bil, med ansiktet nedåt.
Svart man i vit puma tank topp och röda shorts står i dörröppningen av röd byggnad
Två män ler mot varandra.
En liten pojke i randig skjorta fäller stenar för att få vattnet att stänka på honom.
En äldre kvinna gör en formgivning på en vävstol.
En liten flicka leker i en pöl en kall dag.
En hund sätter huvudet på en mans ansikte.
Den lilla flickan sover medan hon kramar sin blå väska.
En flicka som sitter ovanpå en krokodil
Grabben bär en blå jacka och står i grunt strandvatten.
Baby i lekpen med breda ögon
Den tyska herdehunden springer genom snön.
Man sätter upp en bricka i marken.
En vit och brun hund rullar på ryggen i sanden.
En hund skakar av sig vatten
En man spelar en 5-strängad elbasgitarr.
Damen och mannen poserar för en bild.
Byggarbetare lägger stenblock till toppen av en struktur.
Två tjejer går på gatan i shorts och tröja.
Många människor samlas utomhus på natten och äter mat, med massor av ljus.
Ett litet barn som kikar in i en främre torktumlare.
En man i svart skjorta sitter bredvid en gammal kvinna i rosa skjorta på ett tåg.
Mannen i rött pannband klättrar på en sten
Man läser en bok i en frisörbutik på natten.
Två svarta killar, som är på rivaliserande lag spelar basket.
En ung man gör ett förvånad ansikte när han vänder sig till kameramannen utanför sitt kök.
Två män står tillsammans medan en tittar genom kikaren.
Äldre människor sitter tillsammans vid bord och pratar.
En person poserar i snön.
En ensam person som står på några klippor med stora snöiga berg i bakgrunden.
En man höjer armarna på stenig strand.
En manlig vandrare som bär en grön jacka poserar bredvid en stor glaciär.
Någon stirrar ner på en röra på marken.
Den lilla flickan står på en scen klädd som en rosa älva.
En gammal kvinna som fotograferar på en utomhusfotografering.
En flinande flicka sitter i en rosa hjulvagn som glider nerför en grön ramp.
Far och son ler i sängen.
Fem män står i kö framför en röd gardin.
En kvinnlig tennisspelare står redo.
En vandrare står framför berget och håller två käppar.
En brun hund går nära en grön skåpbil och lite skräp.
En svart och grå katt står på en conccption medan två stora hundar stirrar på den.
En äldre kvinna lagar mat i köket.
Två barn, en i röd rock, en i blå rock, sitter vid en sjö.
En fotbollstränare pratar med sitt lag på en fotbollsplan.
En man i solbränd skjorta och bruna byxor tittar nerför fairwayen på golfbollen han just slog.
En kvinna målar tånaglarna när hon sitter på golvet.
En liten hund springer från smutsen ut på gatan
Tre hanar på kanten av vattnet med fiskeredskap.
En elev hoppar upp för att sparka sina klackar tillsammans utanför en skolbyggnad i vintersnöen.
Två hundar dricker vatten i en sjö.
En man med glasögon och en grön skjorta håller fast på väggen.
En kvinna i orange arbetar bredvid en vävstol.
Ett litet barn hoppar på en färgglad leksak på gatan.
En skidåkare fångar luft över snön.
En vit hund leker ute på en inhägnad gård medan det snöar.
En person som har en "fri kram" skylt, kramar en annan person.
En baseball hämtas från en åtgärd som vidtas på ett behandlat fält bevakas av andra.
En kille står och tittar på en annan kille i luften.
Ett litet barn i en röd rock pekar på en handväska i ett skyltfönster.
Ett litet barn står vid kanten av skogen.
En svart hund som hoppar från en flodbank nära ett skogsområde.
Killen som dricker dryck utanför ljust upplyst källare.
Fem asiatiska flickor är på väg på en bana som förbereder sig för att springa.
Fyra män pekar på en mätpinne medan de hukar sig.
Två unga skolungdomar springer för att avsluta sitt lopp.
Tre asiatiska män springer och vinner ett lopp.
Grupp av asiatiska barn klädda i vit polos och marinblå byxor.
En pojke är omgiven av duvor.
En grupp i uniform marscherar med röda skyltar med kinesiska bokstäver på dem.
En kvinna på en skidbacke.
Ett barn som bär en grön tank topp med nummer fyra på det deltar i ett lopp.
Barn passerar en stafettpinnen under en reläkörning.
Det blå laget passerar stafettpinnen i ett relälopp.
Två personer står på stranden och tittar åt höger.
En tatuerad kvinna i svart klänning dricker medan hon sitter vid ett bord i ett svagt upplyst rum.
En man som poserar för sitt foto på en stenig strand.
Toddler stod nära en stolpe med en orange flytväst vid fötterna.
Tre pojkar tävlar mot varandra.
Två tjejer tävlar i en tävling.
Orange hund hoppar över randiga inlägg på kursen.
Två personer som bär svart sitter på en bänk och tittar ner.
En parad av människor i rosa marscher på.
Utanför asiatisk festival med vita ord på röda fanor, en scen av domare bakom en rad röda blommor med massor av asiater stående.
Flera barn på en asiatisk mässa verkar vara engagerade i ett spel.
Barn som håller främmande fanor stående framför en äldre man och kvinna.
En äldre man sitter på en utsmyckad stol med ett bord framför sig.
Två män i en grupp på 4 personer tittar upp på en stor tvålbubbla.
En publik njuter av en utomhusfestival.
Två äldre kvinnor, båda i långärmade jackor med vitt hår, håller händerna nära väggen med graffiti.
Två flickor och tre pojkar sitter på en bänk och skrattar.
Den vita hunden vadar i dammen uppe på berget.
En liten pojke som tittar på en röd vägg
Asiatiska kvinnor som står framför en vattenförekomst och omges av träd med röda löv.
En asiatisk pojke lutar sig mot en stolpe.
En ballerinalärare visar en ung flicka hur hon ska positionera sig.
En pojke läser vid ett skrivbord framför stängda persienner.
Folk går nerför gatan förbi en Lounge &amp; Grill.
Två unga barn är i en hydda.
Ungdomar använder datorer bredvid varandra.
Tre män i en rustik stuga som arbetar med bärbara datorer.
En liten pojke leker på ett djungelgym med ett blått tak och en gul tunnel.
Människan sträcker sig efter något i en plastbehållare utanför.
En vit hund leker med en brun hund på mattan.
En pojke som leker i vatten.
En äldre man i solbränna går över en gata.
En familj går längs en naturstig och skjuter ett litet barn i en röd barnvagn.
En ung pojke håller upp en krokodil till kameran.
Två kvinnor står vid en dörr bakom en annan person som sitter i en röd stol.
Folk shoppar på en marknad med massor av frukter.
En pojke står nära vatten med en sten i handen.
En ung pojke kastade en sten i en damm framför en stor byggnad.
En gammal man spelar gitarr framför en röd hink fylld med pengar.
En sittande, äldre kvinna som fullbordar en målning av en grupp afrikanska kvinnor.
En kvinna klättrar upp för en brant klippa.
En svart hund springer genom ett träskliknande område.
En man och en del cyklar står framför en stor byggnad.
En man som bär en gräs kjol, står i gräset bland en grupp grisar på ryggen nära kusten.
En person som klättrar upp för ett snöigt berg.
En kvinna som bär slöja sitter framför en filt.
En äldre man som sitter framför en bil.
En vit hund med bruna fläckar hoppar genom luften.
En grupp kvinnliga dansare dansar på en scen.
En brun hund med röd väst springer i gräset.
En rodeoman rotar en kalv under en tävling.
Silhuetten av tre män är antingen stående eller sitter i en båt till havs när solen går ner.
En man sitter på en röd soffa bredvid en katt.
Tre barn i baddräkt leker i skum
En man som reparerar en trottoar på en brant kulle.
En man som kastar eller hämtar en lina kastad i vattnet vid en stor båts brygga.
En lerig jeep som kör genom skogen.
En man går mot ett garage, på en dåligt upplyst väg.
En mor och dotter som står framför en graffititäckt vägg.
En fluffig vit hund tittar nerför en brant, gräsbevuxen vall.
En stor båt kör genom hamnen.
Två barn sover i stökiga fåtöljer framför CD-hyllorna.
En falk sitter på en flickas vänstra arm när en man hjälper henne och talar in i en mikrofon.
Två fotbollslag konvergera på målet och målvakten når för bollen.
Barnet i den röda jackan och orange vantar sitter i snön bredvid en spade.
En grupp människor sätter sig vid ett bord för en måltid.
En kvinna som sitter vid sidan av reden och säljer bananer.
2 män sitter ner och ritar på vardera sidan av en staffl i ett rum med en julgran.
Det finns människor som matar får och en hund föder upp dem.
Fem kvinnor i identiska baddräkter håller i ett rep nära havet.
En brun hund sitter framför en kanot.
En brun och svart hund hoppar genom det nyklippta gräset.
En gammal man som bär glasögon ber med sina pärlor när han sitter ner.
Människor som hänger på stranden i baddräkter och avkopplande kläder.
En familj i flera generationer som äter på en restaurang.
Det finns flera kvinnor, vissa bär t-shirts med HSBC på dem, vid en matbuffé.
Ung flicka kramar sin röda nallebjörn.
Flera barn i ljusa färger spelar ett spel av musikaliska stolar.
En trevlig kvartersgata i de vackra gröna kullarna.
Vit fluffig hund hänger ut genom fönstret i en turkos byggnad.
Hunden springer i gräset bredvid vattnet.
En blond hund med floppiga öron springer mot kameran.
En man som håller i en plastpåse står i en dörröppning.
Fyra personer står nära en blå gaffellift.
Ett brunt hår krossas av vinden.
En man med randig skjorta står på scen bredvid en annan person med gitarr.
En fotbollsspelare klädd i blått med en fotbollsboll som förbereder sig för att kasta den.
En man som bär glasögon spelar ett stort mässingsinstrument
En liten flicka tittar ut från en vävd korg.
Duva stirrar på en kvinna i svarta stövlar som sitter på en parkbänk och läser ett papper.
En liten flicka sopar en uteplats med en kvast som är större än hon är.
Mannen som står på bjälken bär en vit hatt.
Stadsartist, manlig, klädd i svart med cowboyhatt som spelar gitarr.
Byggarbetare på en balk som hjälper kranen att placera en annan balk i rätt position.
Man i blå tröja som mäter böjd bräda.
En man som går på sidogatan med huvudet nedåt.
Man på en strand med en baby
En leende man med kort brunt hår i svart skjorta med en öppen orange skokartong.
En dam tar hand om sitt barn.
Två män spelar ut en scen framför en liten grupp vänner.
En kvinna bär en egytisk huvudbonad.
Två unga flickor och en gammal man med grått hår och skägg öppnar julklappar.
Äldre kvinna i rött sötare öppnar en present.
En brun hund ligger på rygg på en vit matta med en grön boll på sig.
En person tittar på en målning medan en annan håller upp handen.
En hummer kör genom en lerpöl flera meter djupt.
En kvinna i svart skjorta kramar en katt.
Damen är vit och säljer saker på gatan.
En hund och en ko står på en bergssluttning.
Två unga pojkar simmar i en pool med grönt vatten.
Två män stirrar på ett flytande föremål.
En kvinna med fötterna på sätena i en tunnelbanebil.
Män som leker med en röd ring ute på fältet.
En pojke som springer på en strand och tittar ut över en stad.
En man i svart shorts glider på en presenning.
En ung pojke i baddräkt och sandaler står i en dörröppning.
Två barn är ute i en liten båt i havet med en större båt i bakgrunden.
Folk går längs trottoarerna i en ljust upplyst stad.
En grupp människor spelar instrument.
En asiatisk kvinna i svartvit tryckt skjorta sitter vid sidan av en byggnad.
En grupp män klädda i tomten klädda spelar musik i ett gathörn.
En tjej som bär en blacker top äter tårta vid ett bord.
Byggarbetare som lutar sig mot under ett tvärgående ljus.
En person är en röd hatt och vinterjacka tittar i fjärran.
En man av afrikansk härkomst står ovanpå en stråle.
En skara ungdomar i förorterna väntar på att en föreställning skall börja.
En person står på en stege och hänger tapeter.
Några personer parkerar sin båt vid en brygga.
Man sitter i en restaurang vid ett bord.
En kvinna i en orange tröja håller i en fotboll och jagas av en kvinna i en blå t-shirt på ett fält.
En man med ryggsäck på att filma något.
En svart och vit hund i en rutig rock bär en mycket lång pinne.
En leende man som står på två skotrar.
En vit hund är luftburen samtidigt fånga en grön leksak.
En person med skateboard sitter på en bänk.
Mannen i blått slår mannen med de röda handskarna medan han blockerar ansiktet.
En man i vit skjorta som äter grönsaker.
En kvinna som håller i en handväska går framför två dörrar.
Ett litet barn som smet nerför en snöig kulle med en blå hjälm
En man spelar akustisk gitarr för en publik inne i ett stort gult och vitt tält.
Fyra Walmart-shoppare i en djup diskussion i livsmedelsavdelningen.
Två personer som bär ryggsäckar och en kvinna i röda shorts står på några stora klippformationer.
Vandrare som går upp för den röda lervägen.
Ett band som uppträder framför en grupp fans.
Ett band som spelar på en ganska liten plats.
En liten pojke äter något och har det över hela munnen.
Band som uppträder på en show.
Två män sjunger framför en liten grupp män med mössor.
En munk visar besökare en av sina ägodelar.
En man i underkläder poserar för en bild med två kvinnor på Time's Square.
Vissa män står vid sidan av motorvägen.
En person med röd hatt står i en snöhög på sidan av en väg medan trafiken går förbi.
En vandrare i en röd mössa som går längs en bergsstig.
En man i blå jacka står på en grusväg i en skog full av träd och ormbunkar.
En hund som sitter i is och snö.
En varmklädd pojke som låtsas att en istapp är en pistol.
En ung man har somnat utanför medan han vilar huvudet på ryggsäcken.
Ett ungt barn med snö i ansiktet kommer ur en blå släde.
En äldre man med glasögon som pratar i telefon.
Två män, en klädd i rött, vitt och blått och den andra klädd i mörk rock, går nerför en kullerstensgata.
Två män i svarta jackor går nerför gatan.
Barn i orange jacka och en hjälm som leker i snön.
En pojke dyker ner i en pool nära en vattenrutschbana.
En grupp människor står på trappan till ett gammalt hus.
En excentriskt klädd man och hans hund sitter på en bänk med gitarr och munspel.
En man som spelar trumpet längs sidan en kvinna som spelar saxofon står utanför i rosa hattar.
Den här kvinnan ligger på betong.
En man med en röd tröja med en pappersbricka som tittar ner på något.
Fyra personer är på en brygga och två av dem sitter på räcken.
En pojke hoppar i en pool medan livräddare tittar på.
En stor grupp människor med broschyrer sitter i en hörsal.
En man med gitarr och cowboyhatt uppträder framför en mikrofon.
Två lantmusiker stör det.
En man på en biltomt håller en pop och väntar på kunder.
Två män jobbar på en cykel i ett garage.
En kvinna och ett barn är utanför en Mcdonald's och det finns en man som sitter inne med en drink.
En man ser ett litet barn måla med sina kritor.
En liten flicka i röd skjorta som spelar på ett djungelgym.
Barnet håller i en tomtefigur.
Fem barn, två pojkar och tre flickor, med flickorna klädda i vita halsdukar, sitter på trottoaren utanför framför ett stort fönster.
Julen på ett torg fullt av folk.
En kvinna i grön väst lutar sig tillbaka med slutna ögon och munnen öppen.
Ett litet barn gråter när mannen i den vita skjortan håller fast honom.
En vuxen håller upp ett barn som försöker åka skridskor.
En man sitter på en vit gräsmatta framför en blå byggnad.
Två hundar, en brun, den andra svart och vit, leker på en trottoar.
En pojke tittar på en ny leksak under julen
Fyra män går nerför gatan i alla svarta dräkter.
Ett barn med en gul ballong går genom en mässa.
En man öppnar en present och poserar med den för en bild.
Människan öppnar presenten av ölflaska kudde.
En tjurryttare försöker stanna på en tjur på en rodeo.
Pojken hoppar ner i en sjö.
En ung kvinna i en muffinsskjorta packar upp en present.
En flicka går bredvid en pool.
En ung kvinna i hatt poserar med en tupp.
Två unga flickor njuter av sin dag i parken med bubblor.
Det finns en person som sitter på en uppblåsbar float i hög snö.
En person i en blå jacka står längs sidolådor och kölar på en livlig asiatisk gata.
En gammal dam bär förkläde i sitt kök, ler medan sked soppa till en annan kastrull.
En tjej i blå baddräkt går över stranden.
En kvinna ligger på magen på en vit kudde och gråter.
En liten pojke kastar snö utanför.
En man som bär svart hatt och rock gör ett ansikte med en folkmassa bakom sig.
Familjens blickar när nyfödda sover i moderns knä.
Det är jul och det snöar också och det är en person som hoppar på en stolpe.
En kvinna och en flicka rider en släde nerför en kulle ståendes upp.
En svart hund bär en orange boll, går på marken täckt av löv.
En ung pojke och flicka som spelar Pokemon.
En äldre person som står i vattnet och håller fast vid en träpåle.
En äldre man och kvinna har monopol på barn.
Två äldre barn håller händerna på ett yngre barn i glasögon medan de hoppar i en bassäng.
En kvinna och ett barn står bredvid en kritbräda på en staffli.
En man spelar akustisk gitarr på en tunnelbaneplattform.
En ung pojke skriver på en krittavla.
En liten flicka färglägger noggrant bilderna av en färgbok.
En liten flicka har en penna som sticker ut ur näsan.
En kvinna i brudklänning går in med en man i kjol.
Två äldre kvinnor lagar middag.
En kvinna i blå klänning som dansar inför en publik.
En manlig bebis färgar en bild med en grön krita och en svagt upplyst restaurang.
Barnet bär en haklapp och sitter i en vuxen'
Tre lättklädda män på en gård ler.
En gyllene hund hoppar i ett försök att fånga en boll.
Hundhoppning ser upp och liten vit boll i luften passerar förbi
En man med glasögon ersätter ett urbatteri medan en annan man tittar på honom.
En ung kvinna och några vänner på en fest.
En man som sitter vid ett matbord och bär en randig skjorta äter en sallad och dricker ett glas rött vin.
En kvinna i gul kostym som ler.
En kvinna läser ett papper högt när en man står bakom henne.
Två män poserar för en bild medan de dricker öl.
En man med glasögon som håller pojken upp och ner ute på en stenfylld gård.
Folk på jobbet i loungen.
Ett gäng killar som tittar på något på en datorskärm.
En grupp brandmän samlas på gatan.
En kvinna med bagage går längs en gata framför en stor annons.
En man håller en hund och en öl medan han sitter i en blommig fåtölj.
En kvinna i pyjamas och en man som ler i en hall.
Vissa kvinnor sätter ljus på en tårta gjord av Marshmallow Peeps.
Två barn tittar genom ett fönster med en vuxen i ryggen.
En kvinna på en restaurang som äter en maträtt.
En polisman pratar med föraren av den blekgula bilen medan tre andra poliser står i närheten.
En ung pojke i en tandläkarundersökning.
Skolungdomar trängs runt ett lägenhetsbord och äter med pappersplåtar och muggar.
En person ger ett rosa pip till en annan person.
Två vita hundar går genom djup vit snö.
En svarthårig man som står bredvid ett podi av trä och plast.
En grupp människor tycker om sitt sällskap med sprit.
En hund hoppar från en brygga och ner i vattnet.
När en åskådare tittar, hoppar en man över en vattensamling som ligger på ett fält av dött gräs, med döda träd i bakgrunden.
En man med hatt kör bil.
En kvinna med en vit tröja kontrollerar blodtrycket på en man i gul skjorta.
En grupp på sex vänner kopplar av i matsalen.
En ung pojke i t-shirt och jeans går på ett gräsfält.
En pojke i blå skjorta får brottas med en rodeo clown i bakgrunden.
Arbetare klädda i jackor och vita hjälmar som går in på en arbetsplats.
Vit fluffig hund kysser får genom ett staket.
Professorn läser namnen på de studenter som har klarat provet.
En ung dansare poserar på ett öppet fält.
En kvinna i vit klänning dansar på stranden.
En surfare som rider en våg i havet.
Ett diagram med en hand visas på en vägg, bakom vilken en kvinna studerar.
En kvinna tittar ut genom fönstret upp mot himlen.
En grupp människor sitter runt ett bord och höjer sina glasögon.
Två personer befinner sig i en kanot på en flod under dimmiga förhållanden.
En äldre kvinna med latexhandskar och man som håller en plastpåse på en fiskmarknad i ett främmande land.
En längdskidare med ryggsäck över en snötäckt bergssluttning.
Flickan i rosa med det ovanliga håret och makeup står vår på den trånga rulltrappan.
Två flickor med hattar springer genom snödrivor utanför.
Fyra personer sitter runt en köksdisk medan man dricker ur ett glas.
Kvinnor står framför en bankomat på ett kasino.
En kvinna i vit skjorta sitter framför en spelmaskin.
Fotbollsspelare skakar varandras händer på fotbollsplanen.
En domare pratar med ett par fotbollsspelare i röda tröjor.
Många män spelar fotboll, medan en publik tittar på.
En ung pojke som stod i ett förfallet skolrum med kritbrädan och ett trasigt skrivbord i bakgrunden.
Mannen i arbetskläder driver en roterande trumma.
En kvinna i maroon springer av andra människor klädda i löparkläder
Två män tittar på andra på stranden.
Två fotbollslag gör sig redo för straff efter en målvakt dra i en match i London, England.
Två fotbollsspelare går på fotbollsplanen.
En flicka med rosa rock och röd hatt går nerför en grusväg.
Står bredvid ett staket, folk samlas för att titta ut mot vattnet nedanför.
En svart hund försöker springa med benen begravda i snön.
En person i svart jacka är snowboard på kvällen.
En gammal man som släpar sina varor i en trehjuling
Två kvinnor som bär traditionell afrikansk dräkt som passerar framför en nedsliten byggnad.
Tre hundar springer över snön med ett däckspår i sig.
Barnen turas om att rida mineraturponny med en vuxen övervakare.
En liten flicka som bär en vit skjorta lägger handen i en fontäns vatten.
Blondhårig man tittar rakt på kameran medan arbetskamraten gör mat.
En man sitter i en båt på stranden med sjön i bakgrunden.
Bricklager som bygger en vägg.
En man i svart hatt och svart rock står bredvid en kvinna som bär en blå halsduk.
2 små flickor gjorde papper platta snögubbar.
En man och en kvinna sitter på en gul soffa och skrattar under en gul tröstare med vita tusenskönor.
Tre barn leker i en vattenfontän.
En kvinna klädd i vitt med hjälp av ett rep för att dra en svart snidad träbjörn på en vagn.
Ett vackert fotografi av en kyrka vid solnedgången med fåglar flyger över och orange-röd himmel
En pojke och en flicka studsar på en boll
En skidåkare ute njuter av backarna på en skarp, cool dag.
En cykel sitter på toppen en uppgång med berg i bakgrunden.
En liten pojke som använder en blå toalett.
Två barn, en i rött, en i svart, glider ner för en snötäckt kulle när de skrattar.
Två arbetare i gula västar försöker fixa något.
En asiatisk man som har tjocka vita handskar, pratar på en mobiltelefon och jobbar på något.
Två män rider scooters genom ett rum.
Det finns två personer, en man och en kvinna, som sitter på en buss.
Barn hoppar och leker i ett hopphus.
Person som håller en frisbee med en vit hund hoppar för det på en väg.
Folk försökte testa ny teknik.
En man sitter på huk nära en brand och håller in något i den.
En kvinna står bakom en utegrill med en blå korg med mat i händerna.
Två vita hundar springer på gräset.
Blå tävlingsbil rider på grusväg med åskådare.
En man som cyklar nerför gatan drar en stor bunt i en vagn bakom sig.
En man och en kvinna pratar med varandra.
En livsmedelsbutikstjänsteman kollar att det är en kvinna med en skadad hand som köper matvaror.
En man i en röd luva som ligger ner i gräset.
En person i snöjacka skyfflar snö.
Olika personer i baddräkter och shorts klättrar stora klippor nära vattnet.
En liten pojke med en brandman hatt på med hjälp av en såg för att skära stjälken av en blomma.
Lokala bybor förbereder sig för en fisketur på denna underbara fiskebåt.
Fyra skjortlösa män, hårt arbetande, på en ställning.
Barn som bär brandmanshatt sitter på marken bredvid en man som håller en handsåg.
Det finns en man med glasögon och en hatt med en svart kostymjacka inomhus.
Damen går förbi en man på en bänk som tittar på henne.
Två män i hårda hattar inuti en struktur tittar på en gul traktor.
En leende arbetare, i en cowboyhatt, som gör murare.
En kvinna i gul bikini topp och solglasögon i en massa människor på en strandpromenad.
Kvinna klädd i rött stående framför flygvapnet män stående i bakgrunden.
En man står framför en fallen byggnad.
Folk är klädda i kostymer på en strandpromenad.
En pojke lutar sig mot en stol medan en annan pojke drar runt honom med ett rep.
En liten flicka i blå klänning som rider på en röd leksakstraktor.
Den bruna hunden springer genom snön
Lokala bybor som åker hem efter en dags skörd.
Ett barn tittar genom persienner på en lastbil utanför.
En pojke gör en kanonkula i en pool medan en flicka tittar.
Ett brunt djur vinkar i ansiktet av en brun och vit tjur.
Ett litet barn tittar genom myntdrivna kikare bredvid en vattenförekomst.
Detta är ett barn i en snöig landskapsspann nerför en kulle.
Två hundar som leker keep-away med röd leksak på blå sträng.
En röd-tjusig, vitskäggig man ler när han står på ett arrangemang av färgglada arrangemang av korgar och dekorationer.
Tre barn leker i en sprinklerpark.
En pojke som bär en röd skjorta dumpar vatten ur en gul hink på en flickas huvud.
Två kvinnor i svarta jackor läser en tidning och ler.
En grupp vänner gör sig redo att åka skidor.
Folk åker skidor nerför ett snötäckt berg.
En pojkes snöslang på ett grönt, blått och gulfärgat rör.
Fem personer håller i instrument och övar musik tillsammans bredvid en byggnad.
Här är en bild av en man pole dans framför sina vänner på en hus fest.
En brun hund och två vita hundar är bundna efter en boll.
Tre personer tar en lift upp för berget i skidorten Adirondack express.
En liten flicka i blå rutor dansar på gräset.
En ung man med en huva stående i ett träskområde med en kamera.
Två ungdomar tar sig genom skogen.
En extrem cyklist, som bär en röd och vit jacka, flyger genom luften på en röd cykel.
En flintskallig, äldre man som leker med en hund.
En ung blond pojke äter en banan medan en äldre kvinna i bakgrunden klockor.
Två unga flickor ska bada nära bergen täckta av snö.
Två kvinnor i medicinsk mask som arbetar i en matfabrik.
Person som dansar på havet.
Två blonda kvinnor poserar framför kameran med en stor grön leksak.
En man och en kvinna skrattar tillsammans.
Ett spädbarn som sover i barnsängen i pyjamas.
Ett barn i en kampsport uniform hoppar i luften med armarna och benen utspridda.
En liten pojke i baddräkt förbereder sig preliminärt för att kliva i den klippiga bäcken.
Folk samlas i en gymnastiksal för en sammankomst.
En brun hund springer nerför en sluttning medan en man följer med honom.
En grupp människor vid ett bord med glas öl leende.
En liten svart hund morrar på en stor brun och vit ko.
En liten flicka med halsband simmar.
Greyhoundhundarna tävlar längs en grusväg med byggnader i närheten.
Tre män står utanför en restaurang och röker och samtalar.
En man slår grillat kycklingben medan en annan kock tittar på.
EN S.C.U.B.A. dykare simmar i djupt blått vatten.
En man ro på sin båt genom mycket stilla vatten.
En liten pojke i röd skjorta som håller en superman producerar och stirrar på en äldre man.
Tre personer går genom en ravin mellan två klippklippor.
Den äldre kvinnan pratar med barnet.
En grupp människor delar en måltid vid ett stort bord på en restaurang.
En brun hund är på väg att hoppa.
En arbetare arbetade aktivt med att svetsa ihop två räcken.
Två män håller ett läkarseminarium, till en liten publik.
En hund simmar i vattnet.
En liten flicka läser en bok i en säng.
Två blonda tjejer äter och en använder ätpinnar.
Skolbarn jagar några duvor.
Ett barn sitter i en stor rund vit stol, läser, nära en rosa bin full av böcker.
Tjejen som äter spaghetti bär en röd jacka.
Den bruna hunden med en röd bandanna sitter med sina tassar uppe på datorn.
En person hukar sig i slutet av en brygga på en sjö.
En mörkhårig man i svart uniform pratar med en man i svart jacka och svart hjälm på en motorcykel.
En man som försöker hoppa i en flotti i vackert vatten.
Några få människor, mestadels flickor, sitter runt ett bord vid en mycket tjusig händelse när de får sina bilder tagna.
En tjej klädd i rosa skjorta, jeans och flip-flops sitter ner och leker med en klubbmaskin.
Tre män som bär gult står bland vägbyggen, en av männen är i ett hål.
En grupp homosexuella män på ett evenemang.
En flicka cyklar på gatan medan hon bär en röd hjälm.
Nygifta par som delar en kyss.
Två män bär gula och orange västar som arbetar vid en avfartsskylt.
Hunden klättrar på uppstoppade djur inomhus, bakgrunds-TV visar brytande nyheter.
Vit man med amerikansk flagga cape och glasögon står i en grupp människor
En man i en tröja som äter en smörgås.
En man som står i kostym och bär glasögon medan han håller ett papper inne i ett tält.
Vägarbetarna kollar vägarbetet.
En ung kvinna i en vit Dior t-shirt lyfter en silverlåda i ett kök.
En kvinna balanserar flera saker på huvudet som är i påsar.
En grupp barn som bär falska näsor utgör en kamerabild.
En ung flicka i grönt leker utomhus.
En grupp barn sitter tillsammans och arbetar med konst och hantverk.
Mannen i gul skjorta och jeans ligger på trottoaren.
En publik som njuter av ett musikband utomhus en vacker dag.
Flera människor väntar på att få spela musikinstrument
En ung flicka klädd i lila läder, övar på en balansstråle i gymnastiken.
Ett litet barn gråter i sina mammors armar.
En utsikt från ett bord med en ung pojke som låg i en äldre människas knä.
En kvinna föder två barn.
En vit och brun hund fångar en röd boll i munnen.
En man står och tittar på folk på gatan.
En grupp unga flickor springer på ett fält.
En liten pojke i orange hatt som springer.
En hund springer på våt sand när en man i gula byxor går längre tillbaka.
Pojken i den röda skjortan är bredvid en blå vägg.
En person i sarong går mot flera blå utomhusparasoller medan han bär på en solbränd väska.
En hund springer genom skogen nära en stuga.
En svart hund med vita tassar hoppar på höbalar.
En man verkar sova i ett hönslager.
En pojke springer förbi en grupp människor med ballonger i ett lopp.
Utsikt över ett passagerartåg genom några lövlösa trädgrenar.
En pojke och en flicka med en uppstoppad rosa björn går längs trottoaren.
Folk som åker nerför en sluttning.
En ung pojke som bär huva, ler och gömmer sig bakom ett träd.
Man springer efter en frisbee med en annan individ rider grisrygg.
Fotbollsspelare värms upp på planen innan ett spel.
Två barn leker i en flod nära en träbro.
En man och en kvinna som håller varandra i handen hoppar ner i vattnet.
Han leker med den lilla hunden.
En man ser på som en annan man försöker klättra en liten stenblock med sin smuts cykel.
Ett äldre par står vid en köpvagn.
En person täckt delvis med en rosa filt sover som en grå och vit katt sover på golvet i närheten.
Hundar tävlar på racerbanan.
En liten pojke i blå skjorta och grå shorts som springer i en park.
Två systrar på en landsväg som jagar får.
Två damer på en trottoar i en stad och en kollar hennes kamera.
En grupp ungdomar leker i fallande snö.
En ung man som bär en rosa och vit randig skjorta sitter bredvid en ung man som bär en brun skjorta.
Två män sitter på en soffa.
En man med svart hår och en grön skjorta kliar huvudet.
En man spelar tangentbordet och sjunger i en mikrofon medan en ung pojke tittar.
En person som svänger på en gunga
En man med långt hår som cyklar ger fredstecken.
En ung man med dreadlocks hoppar högt i luften nära en vägg.
En pojke bär våtdräkt på stranden.
En grupp män står i kö med sina vapen på sin sida.
Kvinna och man tittar på något roligt på en bärbar skärm.
En grupp mest nakna barn som leker på en bro över lite vatten.
En man som sitter på en båt och bevakas av poliser.
En man sitter och dricker en drink med andra människor i bakgrunden.
En grupp människor korsar en flod
En kvinna vadar genom en pool framför ett vattenfall.
Tre pojkar spelar fotboll i gräset.
En gammal dam med käpp korsar gatan i regnet.
Två personer njuter av en naturskön utsikt från en parkbänk.
En grupp människor hoppar upp i luften med sina armar höga.
En stökig tjej på en klubb.
Ett rödhårigt barn sitter och tittar genom ett räcke vid vattnet medan folk leker på stranden på avstånd.
Två personer arbetar tillsammans och serverar mat på en restaurang.
En ung pojke och flicka leker tillsammans i sanden.
En kvinnlig tennisspelare på en blå bana förbereder sig för att slå bollen.
En tennisspelare i en rosa outfit serverar bollen till sin motståndare.
En kvinna som åker längdskidor, med en brun hund.
Två barn fotograferas när de spelar fotboll på ett fält.
Stugor på vintern omgivna av människor som njuter av det vita pulvret.
Tjejen i den bruna skjortan hänger på en blå stolpe.
Två tjejer på tandemcykel, tittar på väggkonst.
En kvinna som bär ett vitt solskydd spelar tennis.
En man undersöker en cykel under en gårdsförsäljning.
En man i kostym och en officer ler mot kameran.
En ung man med grön skjorta spelar en blå gitarr.
Två hundar leker ute i det snötäckta gräset.
Två äldre män framför en buss.
En man i röd skjorta med solglasögon lutar sig mot väggen
En pojke siktar en pil och båge på ett mål.
En man med svart hatt går längs en väg bredvid en byggnad.
Barnet håller i någons arm.
En man och en kvinna sitter vid ett bord med burkar med öl och cigaretter.
Två män, en som spelar säckpipa och en som justerar säckpipan.
Den stora bruna hunden går genom vattnet i havet.
Kvinnan i en blå regnrock går framför en cementvägg.
Den lilla flickan rider sin röda skoter.
Tennisspelare försöker nå bollen.
En kvinnlig tennisspelare står med fötterna isär på en bana.
En kvinna håller ett barn vid ett fönster.
En man klättrar uppför en brant bergvägg med hjälp av säkerhetsrep.
En man når sin höjd för att hjälpa honom under sin bergsklättring.
En brun hund springer genom en hinderbana.
En ung flicka glider nerför en snöbank.
En man hoppar från en ramp på en snowboard.
En skjortlös man med solglasögon tittar på kameran under en strandfest.
En grupp kvinnor och barn står tillsammans bredvid ett fordon och en flod.
En brun hund med grön krage som håller en käpp i munnen.
En tjej i en blå jacka står framför en tråkig publik medan de tittar på något.
En hund springer över gräsfältet.
En person går med en konstnärlig conption framför Ocean Blue Company.
En DJ står under några ljusa ljus med en annons.
En dam med gröna och vita shorts och topp är på stranden klappar händerna.
En hund leker med en fotboll i snön.
Ett barn i en USA jacka skyfflar snö från trappan framför ett hus.
Ett barn som bär röd randig pyjamas ler.
En kvinna hjälper en pojke att göra apbarerna.
En man spelar gitarr.
En man i skägg och glasögon sjunger med när han spelar sin ukulele.
Åtta personer sitter vid ett bord inomhus för förfriskningar.
Tre tjejer sjunger och en tjej spelar gitarr på en scen framför en liten publik.
Ung blond kvinna med röda pärlor, grå tröja märkt GONTAGA.
En person i säkerhet orange kläder ligger ovanpå ett öppet manhål.
Fotografer tar bilder i en byggnad.
En man med skägg och blå skjorta spelar gitarr.
Pojke med en grön och vit fotbollsuniform som springer genom gräset.
En man som inte bär skjorta borstar tänderna.
En grupp människor sitter ute under en grillfest.
En ung blond kvinna och en man som väntar på att gå över gatan.
Ett barn leker med böcker på golvet.
En skjortlös man rakar sig utanför ett garage medan någon åt sidan håller upp en spegel som han kan se från.
En grupp människor organiserar sina kinesiska lyktor.
Surfaren bär en svart kroppsdräkt medan hon hämtar sin bräda.
Två personer står nära en röd skottkärra.
Flera personer står utanför nära metallföremål inklusive några inlägg.
En kvinna som tittar på dagtid himlen genom ett teleskop som är på ett stativ.
En ung pojke i baddräkt kastar sig ut i luften över vattnet medan en äldre man tittar på.
En gentleman klädd snyggt tittar på något på sitt skrivbord.
En ung flicka som äter en skål flingor ur en stor vit skål.
En man grillar kyckling på en grill.
En svart hund försöker fånga ett kastat föremål som är rött.
En äldre kvinna sveper ut på en solig dag
En tjej i en frillig rosa klänning, som dansar på gräs.
En liten flicka i en mjölig, rosa jacka plockar fram en frukt från ett försäljarbord.
En man som bär förkläde står framför lite mat och håller i en blå behållare.
Unge pojke med gul skjorta hoppar upp på den bruna soffan.
Ett barn som bär glasögon och är inlindat i en handduk gråter framför en pool.
En kvinna med vit handske och flera andra.
En man i keps och blå skjorta låtsas kväva en tjej.
En blond tjej som bär Groucho Marx glasögon.
En vuxen hjälper ett barn att åka skridskor.
Barn i ett omklädningsrum på skolan gör sig redo för en pjäs.
En kvinna med ljusbrunt hår sitter över en man med kort medelbrunt hår.
Ett litet barn hoppar högt ovanför ett sandigt fält.
En person som bär våtdräkt surfar på en vit surfbräda.
Person som cyklar nerför gruskullen i skogsområdet
En liten flicka i pyjamas tar en bild med en kamera
En man som ler och binder och förkläde.
En man kör en vagn med trätunnor tvärs över en tom gata.
En man på en båt som står och paddlar på en flod.
En kvinna spetsar en volleyboll när motståndaren försöker blockera bollen.
En gammal man som spelar fiol bevakas av ett barn.
Brudtärnor i guldklänningar och andra ser på som en man i kostym.
Detta är vår paus snabbt tid och vi poserar för fotot.
En man och en kvinna sitter vid ett bord på en snabbmatsrestaurang.
En äldre kvinna i vit skjorta har en röd väska bakom ett glas.
Den vita hunden sprang över kakelgolvet.
Den hjälmade pojken gör ett stunt på en skateboard.
Två män sitter i en liten båt och sprutar vatten på något.
Två män i shorts och flip-flops går framför Farmer's Market.
En pojke klädd i vinterkläder i en igloo
En flicka klättrar på en sten medan någon filmar henne.
Det blå laget, Mustangs, är på en snabb paus, och hoppas sannolikt att kapitalisera med några poäng.
En svart hund springer över ett fält.
En polis på en vit häst patrullerar stadens gator.
Två kvinnor som bär halsdukar väntar på att få gå över gatan.
En kvinna som bär svart vänder sig till en grupp människor i ett kakelrum.
En kvinna och en ung flicka sitter tillsammans vid ett bord och spelar Monopol.
En dam med långt hår och en hatt går nerför en sluttande trottoar belagd med sten.
Barnet som bär den gröna skjortan är på stranden och pratar med några människor.
En grupp människor går mot vattnet på en strand.
Barn lyssnar på en man i blå skjorta.
En grupp människor tittar på ett fält av grönska.
En liten pojke som försöker borsta en kvinnas hår.
Stora grupper sitter runt som en man i en ljusfärgad polo talar framför en stor träbyggnad.
Musiker samlas i ett klassrum för att spela gitarr och andra instrument.
En pojke med shorts, t-shirt, flip-flops och en baklänges hatt sitter i en fällbar stol och fiskar vid en träpir.
En liten flicka i en rosa kofta hoppar från soffan.
En samling människor runt två långa bord uppsättning med olika färgade skålar och tallrikar.
En kvinna arbetar i ett laboratorium med vetenskaplig utrustning.
Dansare, framför Costa Ricas flagga, avslutar sin föreställning.
En ung flicka med håret stående.
En grupp unga ungdomar från Mellanöstern poserar för bilden
Mannen i glas som bär flanell är i klass, skrivande.
En man som bär bilbälte och solglasögon vilar huvudet i en vinkel inuti ett fordon.
Ung man i vit långärmad skjorta som står framför bergen en molnig dag.
En kvinna som håller och poserar ett spädbarn klädd i en hawaiinskjorta på en skateboard.
En kvinna som pratar med folk som sitter runt henne.
En man med glasögon i svart skjorta som spelar trummor.
En man som spelar en orangefärgad gitarr.
En man i vit skjorta kramar en tjej med blont hår på tunnelbanan.
Saxofonspelaren uppträder i gathörnet.
En grupp människor är utanför och går genom en bygata.
Person som ser ut över havet i vördnad.
En kvinna i röd jacka och orange glasögon joggar.
Väntar på hennes poäng efter hennes mumlande rutin är klar.
Armar av fans lyfts till bandmedlemmar när de spelar gitarrer och sjunger i dåligt ljus.
Fyra män i orange västar arbetar på en väg på natten.
En kvinna och ett barn rider i en park.
Byggarbetare på en byggarbetsplats.
En äldre herre står längs stranden av en enorm sjö med en stadsbild över vattnet.
En kvinna med paraply som följer en bil på en skylt.
En liten pojke i gul skjorta klättrar ut ur en lekplatstunnel i plast.
En man lastar Vons kundvagnar på en lastbil.
Ett barn går på en snöig kulle med armarna ut.
En stor hund står i vattnet.
En dam i svart rock och en grå halsduk bär på shoppingväskor.
En mor sträcker sig ner för sitt barn på en trottoar.
Två poliser i Chicago pratar, medan de tittar på en arbetsplats från ovan.
En man spelar gitarr på Joe's Cafe.
Kvinnor handlar på en utomhusmarknad med apelsiner på displayen.
En liten flicka sitter i en barnstol och ser olycklig ut.
En man som går mot en cykel fastkedjad vid en stolpe framför ett stort fönster tidigt på kvällen.
Kvinnan sopar området framför en affär.
En man driver en maskin som en annan arbetare i en orange väst klockor.
En man med skägg och långt hår spelar gitarr.
En ung pojke som går i parken klädd i mörka kläder och mörk mössa.
Folk sitter vid utomhusborden under en brun markis i en lantlig miljö.
En kvinna som bär en rosa hjälm har en tatuering av en infödd amerikan på axeln.
Byggarbetare arbetar på en gammal byggnad.
Fyra hundar leker med varandra och med käppar.
En asiatisk kvinna poserar på piren nära en båt på vattnet.
En man i blå skjorta tittar på tre lastbilar som sveps bort av översvämningsvatten.
En man som cyklar framför en byggnad.
En svart och brun hund som hoppar i luften nära ett fält.
En man står i butiken Tourist-Info.
Vissa människor i ökendräkt står på och bredvid mattor och tyger.
Svart hund på gården på natten.
En man med mörkblå hatt sitter på marken och lutar sig mot en byggnad.
En svart katt kramar en vit och grå hund.
En man spelar gitarr medan en annan man spelar trummor framför en massa människor.
Barn som bär en röd skjorta sitter på en sten i vattnet.
En grupp människor i silhuett spelar på en strand när surfingen rullar in.
En ung flicka leker i sitt rosa leksakskök.
En välklädd, mörkhårig, mörkhyad ung man med öronknoppar sitter och vilar mot ett träd.
En svart hund jagar en pojke i rött och blått.
Två stora hundar vadar i havet
Mannen på en pir tittar på två hundar som står i grunt vatten.
Två kvinnor i vita huvuddukar läste ett sms framför en upptagen affär.
Två unga män i matchande kläder ler.
En brun och vit hund som springer i ett gräsfält.
En man rör vid en stor metallstruktur.
Unga män viftar flaggor i en folkmassa utanför en glasig byggnad.
En man håller flera Tehelka tidningar om ett mord.
En afroamerikansk man med en väska i en blå telefonkiosk.
En man med ett målat vitt ansikte som visslar.
Mannen i röd skjorta står i kö på en restaurang.
En svart och brun hund som springer på ett fält
En man i svart jacka håller en liten flickas hand medan han går nerför gatan
En kvinna med blå skjorta läser för sin son.
En handikappad person med ett ben som åker skidor nerför ett berg med andra berg i bakgrunden.
Man med rickshaw cykel full av mogna bananer.
En man står på en gata i regnet, han håller i ett paraply.
Folk som jobbar i ett kök och lagar mat.
Två små barn åker skridskor över ishockeypinnarna.
Två surfare går längs en klippvägg för att nå vågorna.
En man i en tropisk miljö som håller en kamera mot sitt ansikte.
En grupp människor som sitter på en soffa, en som håller en katt.
Tre män står utanför och en håller en spade full av smuts.
Tre byggarbetare som jobbar på något.
Två personer hänger på säkerhetsrep över en enorm klippa.
Två kvinnor och en man ler mot kameran.
En man lägger sig på en skogsramp medan en annan håller i en fiskespö.
Två barn leker med varandra utanför.
En grupp människor som bär jackor samlas på trottoaren.
En grupp män planterar ett träd.
En grupp och män och kvinnor planterar ett lövlöst träd.
Två män flyttar smuts runt ett ungt träd.
Två unga kvinnor står utanför en blå dörr och en röker en cigarett.
Hockeyspelare väntar på att börja spela spelet.
En brandman på en stege som fixar en telefonstolpe med lågor i bakgrunden.
Gamla händer arbetar på en uppgift.
En man och kvinna klädda i punkrock kläder ses korsa gatan under dagtid.
En kvinna i gasmask använder en symaskin.
En brun och vit hund går uppför snöiga trappsteg.
Pendlingar på ett tåg som ska till jobbet
En kvinna i lila klänning leker med håret medan hon väntar i en lobby.
Barnet i vattnet hålls upp av en vuxens armar.
En skara människor som står bredvid ett skaldjursstånd.
Ett barn bär jeans och en vit tröja.
En liten flicka i rosa hatt är i en frodig grön fält promenader en oxe.
En man som undersöker något under en förstoringslins.
Ett barn står i snön som håller en delvis formad bit snö.
En ung flicka i en blommig klänning omgiven av vattenmeloner
Grupp av barn och vuxna cyklar på en grusväg i skogen.
En kvinna som bär allt blått träffar en boll väldigt hårt medan du spelar tennis.
Toddler pojken bär flygplanskjorta, i barnvagn med stora pärlor.
En man som arbetar på en ångmaskin med ett vattentorn i bakgrunden.
Ett par sitter för att titta på solnedgången från en bro.
En svartklädd man står ovanför en vit hund.
En ung pojke i blå skjorta släpper sin bowlingboll nerför banan i en bowlinghall.
En ung pojke i pyjamas sover på en soffa.
Två flintskalliga män på en parkbänk med små gula trafikkottar.
En man går sin häst på en kapplöpningsbana.
En ljusbrun hund hoppar över ett hinder som har eld i varje ände.
En hund hoppar genom en svart hulahoop.
En skäggig vit man står i en svart kostym med lila slips.
En skallig man kokar på en spis och kastar en knivhuggen fisk i en kastrull.
En stor brun hund som står på bakbenen bredvid en kvinna.
En man som åker buss passerar en man på trottoaren.
En man i orange väst och en mössa står utanför ett damtoalett.
Två pojkar i löparkläder stretching.
En man i kockuniform lagar mat i ett restaurangkök.
Tre män pratar med varandra och dricker.
En ung judisk pojke sitter i en stol på en fest.
En person hukar sig under ett gult paraply på stranden.
Unga flickor springer iväg i en park.
En grupp kvinnor står utanför och pratar.
En äldre man som bär en brun jacka och en hatt står utanför och sträcker sig i fickan.
Två unga kvinnor läser från ett papper till en mikrofon.
Många människor pratar och äter på ett evenemang under dagen.
En kvinna i ett rött förkläde som lagar mat i köket.
En man och en kvinna visar stöd för Mike Huckabees kampanj när de håller upp en skylt.
En tidig man sätter på sig en snidad trämask.
Ett barn leker med ett långt pärlhalsband på golvet.
En mor och en son sitter tillsammans på en säng.
En man bär en picketskylt som liknar en restaurangmeny, medan en kvinna i en rosa, tryckt tröja ger en överdriven pout.
En kvinna i svart skjorta och röd förkläde lagar mat.
Två kvinnor som bär klänningar står ute på gräset medan en av dem håller i en kopp och tefat.
Två personer klädde upp sig och pratade framför ett bord.
En äldre kvinna och en yngre kvinna hälsar på varandra.
Män och kvinnor utanför håller hand för att bilda cirklar.
En brun hund sitter nära en stor sten.
Två personer njuter av havet medan de är under ett paraply.
En vit man som bär en yarmulke står framför en mikrofon med flera andra män i bakgrunden.
Flera personer väljer mat och ökenföremål från en utomhusbuffé.
Två kvinnor, en i vita solglasögon och en grön kjol, den andra i en längre marin kjol, samtalar med varandra.
En hona står med två män som pratar med dem.
Han är på väg att träffa en tennisboll med 3 sekunder kvar.
En man i glasögon slappnar av med fötterna uppe.
En man och en kvinna är vid ruinerna och läser en guidebok.
Ett barn med två fingrar i näsan, täckt av chokladpudding
En man som bär en svartvit hoppsvit joggar längs en väg.
Två män som arbetar med bärbara datorer framför en utsmyckad öppen spis.
En man som bär träningsoverall står mot en stolpe medan andra sitter och lyssnar på något genom hörlurar.
Många hundar tävlar runt banan.
Ett litet naken svart barn står på stranden med fötterna knappt i vattnet.
En kvinna pratar på sin mobil utanför.
En kvinna på en offentlig plats med en gul tanktopp som håller en flaska vatten över axeln
En vacker solnedgång med tre personer i en båt på sjön.
Mannen klättrar upp för ett brant, snöigt berg.
En grupp bandmedlemmar uppträder på gatorna i ett annat land.
Hundarna leker med en tennisboll på gården.
Trött på att läsa sin bok tar en ung man i randig skjorta en tupplur i biblioteket.
En liten hund på ett kedjat koppel står ensam i en skuggad hall.
Fyra personer är i någon typ av cement byggnad med nummer 93 målade på väggen.
Lille-pojken står bakom en glasdörr med röd hatt och svart jacka med en kvinna som står alldeles utom synhåll på trottoaren.
Cykelförare passerar en utsmyckad byggnad med en klocka.
En man med glasögon och en röd ryggsäck som står framför en tegelvägg
Rida en röd motorcykel, med lämplig utrustning.
Två män samlas i lobbyn i en byggnad.
Två personer går i en öken.
En man sprejar en cementbil med en slang på en trottoarkant när en man går förbi.
En man skyfflar snö framför ett hus.
En äldre man som bär vinterrock och jeans står framför en stor, välvd blomstervagn.
Den unga basketspelaren flyttar in i fronten.
Skakigt klädd kvinna i svart väntar i en restaurang med andra beskyddare.
Damen i rosa går förbi nån som håller i blommor.
Några män sitter på stolar och står under ett stort rött paraply.
En kvinna säljer grönsaker på gatan.
En kille som bär parka går på en tom trottoar.
En flickas fotbollslag går in i en kurragömma.
Två män sågar en trätavla som försöker slutföra sitt projekt, medan en av dessa två män röker en cigarett.
En man bär en bricka med glasögon.
En flintskallig man som springer på ett löpband i vit skjorta och randiga shorts.
En grupp män slipar sten under dåliga förhållanden.
Två män i ett garage lagar motorn till en bil.
En surfare vid en bro i dimma förhållanden
En ung flicka glider nerför en snöslänta i en röd släde.
En lokal konstnär uttrycker sig på en vägg vid sidan av en gata.
En kvinna målar den andras ansikte för en karneval.
En kvinna drar upp en uppblåsbar båt i vattnet.
En kvinna som håller i en vattenflaska springer på stranden.
Många människor av indisk härkomst bär ljusa, färgglada kläder &amp; går upp branta trappor.
En stor svart hund bär en blå boll medan två Corgis springer vid hans sida.
En liten pojke tittar på en slottsvakt utanför en liten svart hydda.
Två hundar leker i den vita snön.
Två medelålders män spelar gitarr på en scen.
En gammal kvinna som går längs en trottoar med byggnader som är fulla av graffiti.
Några barn i vitt och rött spelar fotboll.
En man i ett förkläde står i ett kök och arbetar med en industriell blandningsskål.
En grupp människor är utanför en tegelbyggnad.
En utsikt över ett europeiskt stadslandskap fullt av många förbipasserande.
En pojke med en röd ryggsäck som går längs en stig.
En kvinna med pandamössa och hörlurar står framför en man utanför i snön.
En kille som hoppar framför nån intressant väggkonst.
Ett litet barn skyfflar en snöig uppfart med en ljus orange spade.
En ung man med ett glatt uttryck kastar upp bitar av färgat papper i luften.
En man i rutig skjorta kastar en yxa vid en vägg i sitt garage.
Mannen, sonen och säljaren ler medan de håller souvenirtidningar.
En vacker utsikt över bergen en snöig dag.
En schäfer leker med en röd boll.
En pojke och en flicka klädda i snödräkter, hoppade i luften med händerna upphöjda i massor av snö.
En man beige skjorta som tar en drink.
En ung i en vit klänning som står framför ett stängsel och en fontän.
En man håller en skål bläckfisk.
En slaktare som skär fisk för försäljning på marknaden
Hund travande med en gummianka i munnen
En grupp unga vuxna samlas på golvet för att spela ett komplext brädspel.
Två hundar slåss om en pinne i ett översvämmat fält.
En mamma och son njuter av en dag i parken.
Folk går på gatan.
En sky-vy på en restaurang med utsikt över människorna i båsen.
En pojke matar fåglar i en park.
Två män och två kvinnor står vid fönstret i en biljettbås.
En vacker dag att ligga vid havet och vänta på vågorna.
Fyra cyklister rider längs en grusväg mellan två stängseltrådar.
En ung flicka som övar på sin kastrull.
En man sitter vid våra dörrar bredvid kartonger och spelar ett instrument.
Arbetare som bär hårda hattar och ansiktsmasker bearbetar avfall.
Ett barn i rött hoppar på ett rött föremål medan andra skrattar.
En kvinna läser en bok på en tunnelbanestation.
En kvinna i en röd sport-bra springer på trottoaren förbi ett tegelstängsel.
En tjej med färgat rött hår klädd i randiga kläder som pratar på en mobiltelefon.
En person står mellan två gigantiska statyer som ser ut som ansikten.
En präst gnuggar ett kors på en mans panna.
En man leder en karavan på sex kameler och deras ryttare uppför en sandig kulle, med klippiga berg i bakgrunden.
En äldre människa hukar sig ner och håller i en käpp.
Målare i röd overall målar en stor dörr från blått till grått.
En man som rakar en annan man i en frisöraffär.
En skara unga människor i vinterkläder som väntar på tåget.
Hunden går genom det kalla vattnet.
En vit hund hoppar upp för att fånga en fotboll i anlagda gräsyta.
En man med mörk topp och vita byxor ligger ner i skuggan på parkbänken.
Vuxna i vinterjackor och hattar svingar kvastar på en liten gul boll medan en svart hund tittar på.
Mannen och kvinnan sitter vid ett bord.
Barn spelar basket på en bana.
Flera kvinnor sitter i stolar framför en vägg av speglar.
En husvagn med gröna och röda fordon som går upp för ett berg.
En man klädd i vinterkläder är på stranden med en hund.
Ett litet barn står framför en dator på ett affärskontor.
En skulptör i en blå tröja som skär en bit sten.
En kvinna försöker korsa vägen innan en man på en röd skoter.
En äldre kvinna tittar på en tonårspojke
En stor grupp människor klädda samlas lättvindigt för att dansa.
En äldre man med glasögon fixar en leksaksbrandbil medan en liten flicka leker med den.
En kvinna på en mobiltelefon går uppför trappan i tunnelbanan med en annan passagerare i närheten.
En man som säljer eller köper apelsiner på en vagn i en affär utanför.
En pojke i rött hoppar bakåt på sanden på en lekplats.
En pojke hoppar på de ljusa kuddarna.
En brun hund och en fläckig hund käbblar över en hundleksak.
En man i en tröja som lär sig sticka.
Kvinnliga skylthållare tar skydd under paraplyer under en regnstorm.
En grupp kvinnor sitter runt bordet.
En grupp kvinnor sitter nära varandra och stickar.
Flera kvinnor samtalar runt ett bord.
En vit hund i svart rock står i snön.
En grupp människor besöker i ett mörkt upplyst rum.
Tre honor hänger medan de andra tre honorna går sin väg.
En enda man som dricker en mugg grön vätska
En grupp människor på en fest med två kakor på bordet.
Många gamla kvinnor är scenkonst och hantverk.
En skara människor är på gatorna och en del har facklor.
Ett par människor är klara med att skyffla en stig.
Män som arbetar längs sidan en fisk och chips restaurang med en soptipp lastbil.
En man tittar på sin unga dotters reaktion på en hemgjord födelsedagstårta.
Folk springer och går in och ut ur en liten bondgårdsstad.
En man klädd i svart går på en isig trottoar
En liten flicka i en brun topp och rosa byxor balanserar en skål med växter i det på huvudet.
En grupp människor står på gatan.
En hold man i grön jacka läser en bok längs en grusstig.
En ung pojke som håller en basketboll på väg att skjuta.
Sex små barn i rockar samlas runt en matvagn som säljer kastanjer för 2,00 Euro.
En byggnadsarbetare övervakar någon som gräver med en maskin.
En massa människor sitter på en stadion.
Bilderna dyker inte upp, så jag antar att bilden är underbar.
Två pojkar äter äpplen leker på en cement bil barriär
Pojke med målat ansikte går runt ett spår.
Ett band är på scen och spelar musik, ledd av en man i kostym.
En kvinna ses läsa genom ett tunnelbanefönster.
Unga flicka i rosa klänning leker med pojke och en boll
Flera personer klädda i blått, en snurrar ett band
Två hundar leker med en tennisboll i snö nära ett träd.
En svart man som står ensam ute i en lång överrock.
En flicka ler som en motorcykel med två vuxna och ett barn passerar förbi här bakom.
En ung pojke som tvättar ett fönster.
Kvinna i rosa topp rider en cykel längs sidan en man jogging längs vattnet.
En mamma och ett barn på stranden med segelbåtar i bakgrunden.
En man läser en annons på en busshållplats, medan en annan man sitter på en bänk.
Två pojkscouter fyller hink med vatten från ett handfat
En man klädd i vit skjorta med vita shorts målar en vit vägg svart.
Ett äldre par som njuter av en julmåltid.
Det finns två killar som spelar gitarr hjälte på en offentlig plats.
En liten pojke i en grön tröja som leker med sitt leksakståg.
Kvinnan på gatans fönsterbutiker framför butiken, Louis Vuitton.
Sex personer försöker flytta en bil på en snöig gata.
En man i en blå tröja spelar ett sportspel på Wii!
Två tjejer spelar instrument i en grupp.
En man står på en stor klippas klippkant.
Ser ner på nån som klättrar på en klippa över vatten.
En man som hanterar en guld vas typ objekt med 2 andra tittar på.
En mamma drar sin dotter på en släde i snön.
Tre personer i skidutrustning står bakom en "ingen skidåkning"-skylt.
En liten grupp människor står och pratar med varandra utanför.
En kvinna som bär visir spelar piano utomhus.
En blondhårig pojke tittar på en konstig humanoid robot.
Någon dinglar på ett rep från en klippa över havet.
En bergsklättrare med vit hjälm stöter bort.
En hund som sträcker sig över sandlandskapet framför folk som tittar.
En ung pojke som kissar på sig blå shorts och klumpar som håller i en fotboll som springer från andra pojkar.
Collie står utomhus på ett sandigt område.
En grupp tjejer som hänger på en våt sandstrand.
En ung pojke kastar sin boll i luften utanför.
En ung man ser en liten flicka gå i gräset.
Två delfiner hoppade upp ur vattnet i det här zoot.
En kvinna med röd hatt och svart rock.
Två unga flickor tränar för att hålla jämna steg med att spela fotboll.
Lilla flickan sparkar stenar på stranden med sin hund.
Tre barn hoppar medan en äldre man tittar på från en rad stolar i närheten.
En ung man som plockar på sin gitarr i ett väntrum.
Två peoplw med toppen av huvuden på gräs.
Tre hundar som leker på en gård tillsammans.
Vissa tittar ut genom fönster i en stor byggnad.
En liten pojke i svart surfar.
Två grå hundar springer tillsammans över det gröna gräset.
Den tyska herden går i vattnet.
En ung pojke är på baksidan av en annan person som bär hatt.
En sångare och två gitarrister spelar på en färgglatt upplyst scen.
En äldre gentleman bär en utstuderad huvudbonad som håller en vit hund som har fått sin päls färgad flera färger.
En hund bär en käpp genom skogen.
Två hundar, en stor och en liten, leker tillsammans i gräset.
Fyra personer rider på tunnelbanan.
En skallig man som sitter på en scen och spelar gitarr.
En man i blå och vit skjorta sitter.
En grupp campare äter middag nära sin eld.
Flickan leker tillsammans med bilderna på den stora skärmen.
En brun och svart hund jagar en svart hund i snön.
En rödhårig hane rakar ansiktet.
Flera människor går på en regnig livlig gata i Asien med tydliga paraplyer.
En flicka spelar ett tv-spel på en skärm i naturlig storlek.
En man står framför en byggnad med hjärtformade ballonger och en kvinna går över gatan.
En skjortlös man arbetar på en byggarbetsplats.
En man utan tröja jobbar på sidan av en byggnad.
En fotograf står med en pojke och hans fotoutrustning.
En stor hund springer genom ett fält med en mindre hund.
En man som bär svetshjälm svetsat stål.
En brun och svart hund går i den vita snön.
En kvinna och en liten flicka poserar för en bild med en lama på toppen av en bergssluttning.
En skjortlös, skäggig och mustad man tittar genom ett hems dörr medan en katt sitter på nedre trappsteget av ingången till hemmet.
En åsna som drar en bil med en man på
En blek pojke som leker i en grop av blå bollar.
En utländsk dam som samlar grönsaker.
En hund springer i snön, ett staket i bakgrunden.
En ung pojke som ler och håller i sandaler.
En handskeman går på en trottoar nära en orange skåpbil.
En grupp människor går utanför ett utställningstält.
En kvinna pratar med två poliser i gula jackor vid ett utomhusevenemang.
En snowboardåkare som gör ett trick när han springer.
En man lägger sig för att vila i en träkonstruktion mot en byggnad.
En grön fisk hoppar upp ur vattnet.
En man i svart t-shirt tittar ner när han dricker.
En man som cyklade en dimmig dag.
En kvinna med rosa hatt tittar på en rosa bil med lastbilen öppen.
Kvinnan i blå jacka visar upp sin vintagebil framför Nathalies dockhus.
Två kvinnor i solhatt går arm i arm nerför en stad gata med portmonnäer.
Folk går runt och skrattar utanför.
En kvinna i en grön tank topp med locktång i håret har makeup appliceras på ögonen framför en leopard print bakgrund.
Brunett kvinna fixa blond kvinnas hår.
En kvinna med gult handledskorsage talar till den blonda bruden.
En man i solglasögon sitter med sin flickvän på ett bröllop.
Folk ler medan de står i kostymer och klänningar.
En man och en kvinna ska gifta sig utomhus.
En man och en kvinna gifter sig ute en solig dag.
En brudgummen och bruden tar sig nerför gången som man och hustru.
Män och kvinnor vid en formell funktion när en kvinna i en vit klänning bär en bukett med röda blommor.
En kvinna leder tre små pojkar i fotboll uniformer.
Tre kvinnor i klänningar är utanför och tar emot hors d'oeuvres från en cateringfirma.
En sjaskig hund med en leksak i munnen.
En pojke verkar dansa till musik i en byggnad fylld av människor.
Mamma med barn tittar på blå fisk.
Fyra barn står och poserar för ett foto.
En person använder ett långsökt nät för att fånga något i luften.
En man som bär gröna vattentäter går på en gräsbevuxen klippa och bär på några pingviner.
En man med en kamera studerar sitt arbete.
En ung man i vit skjorta och guld och svart hatt sitter korsbent.
En pojke hänger på remmar på ett tåg.
En ung flicka viker ett vitt klädesplagg från en tvättkorg.
Två personer gör musik med gitarr och tangentbord.
En kvinna som bär en rosa boa cyklar nerför en gångbro.
En ung man som står på brandstege i en stadsbyggnad.
En kvinna i grön skjorta och blå hatt spelar tennis.
En man klädd i blått jonglerar inför en publik.
En kvinna i jeans sover på en man.
En hund som bär jacka, kastar en leksak.
En man håller i skrevet med skjortan upphängd och avslöjar magen, samtidigt som han bär en daggtrasa.
En man som snurrar en skateboard i händerna medan folk tittar.
Barn är mycket glada över att se en papegoja äta mat ur sin hand.
En vit hund plaskar genom vattnet.
Byggarbetare arbetar med en tung maskin bakom en orange och vit randig barriär.
En liten pojke som upptäcker växter som växer i en pöl vatten.
Två lag spelar fotboll, det ena försöker ta itu med det andra.
Asiater äter i en restaurang med orange motiv.
En korthårig man i en mörk kamouflagejacka spelar saxofon i ett gathörn medan folk tittar på i bakgrunden.
Två hundar springer längs en stig full av döda löv.
En liten pojke häller vatten från en hink på en annan liten pojkes huvud.
En vuxen vandrar i snön med ett berg i bakgrunden.
En ung pojke spelar basket i en officiell match.
Tre killar sitter på en bänk utanför en dryckesaffär och pratar.
En stor hund jagar en liten hund på sanden.
En snowboardåkare i vitt svävande genom luften.
Barn, som visas i en flygbild, leker i ett typiskt familjerum.
En kvinna går nerför trottoaren med en plastpåse.
En hund går genom snön i dagsljus.
Två hundar springer över ett gräsfält.
Det finns fem skidåkare, med ryggsäckar, i snön.
En pojke håller en basketboll i en hand.
En snowboardåkare i grå byxor hoppar.
Två bergsbestigare tittar framåt på en snöig stig.
En snowboardåkare lutar sig mot sin snowboard medan han tittar på utsikten över dimmiga berg
Svart hund springer väldigt fort.
En man i en brun jacka som står framför en öppen verandadörr.
Två bruna hundar springer genom ett fält med en röd leksak
En person målar ett foto av en hund, baserat på ett foto av en hund.
Man pratar på mobil utanför en juvelaffär.
En grupp skidåkare går upp för en lutning i snön.
En äldre man står bredvid en yngre man med hörlurar
En skjortlös man med glasögon och vått hår som rakar ansiktshår.
Människan säkrar ett stort betongblock.
En man i grå jacka som sitter på en grön bänk och klappar en svart hund i röd krage.
En man i läder tar en bild av kristall.
Ett äldre barn som ser ett litet barn leka med en lång vår inne i ett hus.
Två små vita hundar som leker
En liten flicka som håller i blommor går bort på en stig en solig dag.
En man arbetar på att bygga ett skyddsrum av stockar och vassrör.
En man, en tonåring och två pojkar blandar en hink med vätska på en gård.
En grupp passagerare umgås medan de väntar på en busshållplats.
En man och kvinna som bär vinterkläder försöker sälja olika föremål på ett bord utanför.
En pojke med orangefärgade stjärnglasögon sitter och håller i en leksakshammare.
Två män utanför tittar på metallföremål.
En pojke kollar ett system på datorn.
Två äldre personer som intervjuas av en kamerastyrka som står nära en grön metallbil.
En hund tittar försiktigt på den bruna hunden som utreder hans område.
En man med svart hatt sitter på en pall framför en grön dörr och bredvid högtalare.
En pojke och flicka plaskar runt i havet.
En man som håller snorklingsutrustning hoppar ner i havets gröna vatten.
En man som står på gatan.
En man lägger sin hand på en annan mans rygg och de är båda på en båt.
Det är en vacker dag för ett utomhusbröllop.
Många människor handlar på en inomhusmarknad.
En ung pojke springer genom bubblor.
Åtta personer njuter av det roliga i flottar och skönheten i ett vattenfall.
Flera människor går nerför en stig.
En man i en blå och lila randig skjorta och hatt går förbi en tegelbyggnad.
I det här fotot säljer en kvinna marknadsföremål.
Det finns en monter under ett stort blått och rött paraply med ett stort sortiment av produkter och det finns flera personer som tittar igenom produkterna.
Ett barn som gör ett sandslott på stranden.
En manlig dirigent som bär alla svarta leder en orkester och kör på en brun scen och spelar och sjunger ett musiknummer.
En ung pojke i en grön hjulpipa med en flicka som knuffade honom.
Killar i en frisersalong en kille som håller upp ett finger.
En lagspelare tar sig tid att kommunicera med media.
En svart och vit hund som bär kragar skakar av sig på dött gräs.
Lilla flicka som ligger i många färgade plastbollar.
En man med skägg sticker ut i färg.
Här är Rod Stewart i Konsertsång Live med Pat Benatar.
Det finns fem sångare på en scen, tre kvinnor och två män.
En hund springer genom det höga gräset.
En kille med solglasögon sitter på en båtfärja i solen.
Hunden går längs en strand vid solnedgången.
Thre är en shot av man med ryggen vänd i en stad.
Två svarta hundar springer på gräs.
Två medelålders män försöker operera vad som ser ut att vara en förstoringslampa av något slag.
Två flickor som målar i en färgbok vid ett bord.
En man i röda badbyxor står i snön på en klippa ovanför vattnet.
En familj står i en snöig skog.
En grupp ungdomar klär sig i ett glest rum.
Två män i vita skjortor och breda vita byxor utför kampsporter.
Två hundar tycker om att leka i snön.
En ung flicka som läser en litterär klassiker "för att döda en hånfågel".
Två kvinnor i en bubbelpool med handdukar på huvudet skrattar.
Skiiers på toppen av ett berg.
En man i en brun rutig skjorta säljer bakverk från en blå varuvagn.
Folk på marknaden plockar ut och tittar på frukt.
En man i blå träningsoverall och en kvinna i brun jacka och bruna stövlar går tillsammans.
En ung man med brunt hår som spelar gitarr.
En grupp män sitter på röda stolar.
En hund bär en tidning genom ett kök.
En man i vit skjorta som visar en ung pojke hur man gör bröd i ett bageri.
En hund går ner för en ramp, tänder bar.
En grupp män sitter runt ett bord som har tomma flaskor på sig.
Två basketspelare tittar på bollen.
En man åker skidor nerför en snöig kulle medan han kastar en lång skugga.
En kille som utför tricks framför barn med coola baseball fladdermöss
En man läser en tidning i en kinesisk mataffär.
En tjej som bär hjälm åker skoter.
En äldre man som arbetar med flera strängar.
En bebis som håller i en skallra ser väldigt ledsen ut.
En pojke surfar mot stranden på en grön surfbräda.
Kvinnan vilar sitt huvud på en böjd kudde.
En ung kvinna bär en brudslöja utanför en kyrka.
En man och en liten flicka i rosa klänning
En man sitter på en bänk med armen runt en dam.
En gyllene hund går försiktigt runt en frusen damm.
En kvinna ler och sätter sina knytnävar i luften i glädje.
En man som bär en blå skjorta som håller i en kedja.
Folk sitter i soffan och skrattar.
En liten pojke hoppar från en stol till en annan.
En hund hoppar upp i luften för att fånga en boll i munnen.
En man med en bock som lutar sig mot en vit skåpbil.
En kvinna med mörkt hår som bär orange bikini lägger sig på en korgstol.
En man i svarta kläder utför ett stunt att svälja tända facklor.
En hund sitter i en bil och tungan sticker ut.
En man som sover ute på marken.
En man i orange arbetar på en byggarbetsplats bredvid en stor lastbil.
Två pojkar åker skridskor med andra människor.
Fem vuxna och ett barn springer mitt emot vågorna på stranden.
En man är upptagen med att putsa en palm.
En man i svart t-shirt tittar på en meny.
En vit hund löper längs en klippig strandlinje.
Mannen står nära tåget vid tågstationen.
Ett skjortlöst barn leker med en rosa ballong på en trottoar.
Man och kvinna dansar tillsammans med pengar över hela golvet.
Saker djur priser människor kan vinna genom att spela en karneval spel.
En kvinna ser det som en spegelreflektion och använder en mascarapenna på sitt vänstra öga.
Ett par beskyddare på en jazzklubb.
En man på en motorcykel som utför ett trick högt i luften.
Pojken kommer nerför kullen i den röda vagnen.
En man med gul skjorta står framför en man som spelar ett musikinstrument.
Två hundar leker i vattnet med en pinne
Ett barn kryper på golvet och tittar på en duva.
Han jobbar hårt på jobbet på gatan.
En person kommer nerför en gul vattenrutschbana i en pool.
Manlig matarbetare grillar kött på en pinne.
Två unga violinister går mot kameran från en dörr.
En grupp människor dansar på en orientalisk restaurang.
Tre män är ute vid solnedgången och gör olika aktiviteter, bland annat hoppar, sitter och leker med en fotbollsboll.
Tjejen träffar volleybollen.
Man i Dr Pepper logo skjorta ligger på en blå filt, med armen runt en leksak tuggande spädbarn.
Två pojkar spelar flaggfotboll.
En man som sover på en annan sovande mans knä på en parkbänk.
En grupp människor som går uppför en gräs kulle.
Person på snöskidor luftburen över snö med grönt träd i bakgrunden.
Tre små barn på trehjulingar tävlar nedförsbacke.
En tandläkare undersöks av en man och en kvinna i blå skrubb.
En ung man som går förbi ett fruktstånd.
En person som bär en tröja med huva och jeans står på ett träd som har fallit över en bäck.
En grupp människor äter tårta på en kontorsfest.
En man är klädd i en svart skjorta samtidigt balansera ett runt föremål på baksidan av sin hand.
Två cowboys tittar i baksätet på lastbilen.
En man är synlig rider en svart häst med en brun häst och tjur i bakgrunden.
Två cowboys från Latinamerika eller Sydamerika rider hästar och jagar en tjur.
Två män på hästar jagar en ko en solig dag.
Barn leker på gården
En man i en roddbåt ro över blått vatten.
En grupp barn leker i ett museum.
En grupp människor rider hästar i gröna västar.
En kvinna som håller tennisracket på en bana.
En man och en kvinna i blå klänning spelar tennis.
En kvinna håller i en tennisracket.
En tennisspelare i röda kläder håller upp sin tennisracket.
Ett barn som ligger mitt i fyllda leksaker och filtar.
En kvinna bär ett barn på ryggen.
Pojken springer över planen med basketbollarna.
Två män båda bär vit t-shirt står bakom disken, båda håller knivar.
Tre brandmän står i en hiss.
En leende, glad-framträdande blond kvinna med ryggsäck stannar för att le mot kameran.
Barnet sitter i en barnstol.
En terrierblandning fångar en frisbee i luften.
Mannen i rocken har guld på skägget.
Ung asiatisk man hoppar upp på toppen av en vadderad rektangulär metall struktur.
En liten pojke leker på en våt stenyta.
Unga kvinnor med gröna mössor som böjer sig ner för att plocka upp en korg från ett fyrabent skrivbord.
En ung asiatisk pojke håller i en liten, vit, långhårig hund.
Vänner och familj dansar på en strand vid sina fordon.
En indisk kvinna poserar för kameran i sina ljusa kläder.
En ljusbrun hund med en mörk krage som sträcker sig genom gräset.
En man i svart skjorta och kamouflagebyxor täckta av grädde.
Fyra män med skägg som står upp och håller vita tallrikar.
En liten flicka sparkar upp i luften.
Vit hund med öppen mun springande i snön.
En asiatisk kvinna och en liten pojke cyklar tillsammans.
En leende indisk kvinna som kör en blå lastbil klädd i en färgglad orange, grön och vit outfit.
Två personer hoppar från en sanddyne på en strand
En man, som bär randig skjorta, driver ett mikroskop i ett laboratorium.
Ett barn sitter i ett hål fyllt med vatten.
Den bruna hunden går längs en gräsbevuxen stig med tungan ut.
En svart hund springer med en vit hund
Två stora hundar springer tillsammans genom gräset.
En hund rullar i gräset.
En pojke i rött förbereder sig för att glida ner för en blå rutschkana.
Flera män på hästryggen stirrar in i en bergsbakgrund
En dam med en fin kostym och huvudbonad medan hon dricker från en burk.
En valp bär en tennisboll i munnen.
En kvinna med fem barn runt omkring sig med ett leende på läpparna.
Människan paddlar en kanot genom stilla sjövatten
En del människor går över en grön bro över en flod.
Två unga män hjälper en annan man i ett butiksrum.
Två pojkar klädda i slitna fasta färger kläder står sida vid sida medan en håller en yxa.
En man som sitter vid ett bord med hjälp av en bärbar dator.
Ett barn vänder sig om med ett föremål i handen medan någon passerar bakom honom.
Två kvinnor samtalar i ett konstgalleri.
En person och deras bruna hund åker en sväng i en roddbåt.
En brun hund som sitter på gräs
En vit hund springer med ett orange staket bakom sig.
En man och en pojke tittar in i ett tält med en blå filt i.
En kvinna med tennisracket på väg att svinga mot en boll.
Kvinna i vit skjorta och svart kjol spelar tennis.
En kvinna med en huva i tröja och svarta byxor med en hästsvans som spelar tennis.
En blond hund som leker med en färgglad hundleksak.
Två tjejer med långt hår står framför ett rörigt bord.
En tennisspelare höjer sitt racket för att slå bollen.
En liten flicka går på en stig i en inomhusträdgård.
En kvinnlig tennisspelare som ska slå bollen.
En brunhårig kvinna i en beige jacka skriver på ett papper på ett rosa bord.
En kvinna med vit kjol spelar tennis.
En blond kvinna som spelar tennis, framför en blå reklambakgrund.
En indisk man och kvinna sover på kollektivtrafiken.
Ett barn som ler när de kastas i luften av en vuxen.
En kvinna med grönt hår svingar mot en pinata.
En svart och vit hund springer över snön vid ett träd och en bänk.
En tennisspelare som samlar tennisbollar i en tennisbana.
Kvinnor på tennisbana står framför nätet och håller i en bok.
En glad tennisspelare i en vit sportbehå.
En tjej med vit topp och gula shorts spelar tennis.
Det finns en kvinna i gult spelande tennis.
En ung tennisspelare sträcker sig för en boll på en lerbana.
En kvinna i en vit tennis outfit som spelar tennis.
En kvinna i en blå sport outfit är på väg att slå en tennisboll.
En man som går framför graffiti en molnig dag.
En äldre och yngre kvinna, både med tenniskläder och racketar, ler sida vid sida för kameran.
Barnen gör snöänglar bredvid varandra.
En kyrkogårdsarbetare gräver, eller fyller en grav, en annan person är på sin mobiltelefon, lutande på en gravsten.
En person i pälskrage går förbi en staty.
En man och en kvinna använder en maskin inbyggd i väggen.
En afroamerikan som går nerför gatan i en ljusfärgad skjorta.
En pojke klädd som en cowboy klappar ett fyrbent djur med horn och en sadel.
En ung cowboy fascineras av en kamels närvaro.
Tre barfota barn roar sig och ler i en inomhusmiljö.
En man med muskulösa armar utför gymnastik.
En man i rött tights balanserar på en bjälke med benen i luften.
En kille kommunicerar med någon i en bil.
Honan är redo att slåss om det behövs. Hon är tränad.
Den svarta och vita hunden hoppar för att fånga en leksak.
Två små barn knuffas på en däcksvinge med snö på marken.
En äldre kvinna som deltar i en ceremoni.
Stor brun hund hoppar över en buske i ett gräsbevuxen område.
En gymnast hänger upprätt i ringar.
En svart pälshund hoppar i luften bredvid en annan hund.
Två unga pojkar som ser sin far använda en stand up mixer.
En brun hund leker med en röd hund i snö.
En liten blond tjej på en klättervägg.
En man har sina skor lyste på trottoaren på gatan fodrade med parkerade motorcyklar.
En man kysser en kvinna på kinden.
Tre barn och en vuxen som går på en stig.
Flera personer sitter på en bänk före solnedgången.
En man röker en cigarett och den andre möter sin blick.
En hund som simmar med en käpp i munnen.
En man som bär stora snöskor springer in i en till synes fullsatt skidort.
En gråhårig man sitter utanför och pratar i telefon.
Två små barn kurar runt en kvinna på gatan mellan två gröna och gula vagnar.
Två män sitter och dricker.
En brun hund leker med en röd leksak medan en annan brun hund går mot kameran.
En kvinna glider bakåt i snön.
En man som bär t-shirt och blå jeans hoppar från en klippa vid en stor kanjon.
En man och ett barn sparkar en gul boll i ett öppet fält.
En pojke i blå skjorta hoppar ner för trapporna på en skateboard.
En bowlare kastar en boll längs banan och försöker träffa två stift.
En kvinna i rosa hatt hjälper en liten flicka i vit hatt med sina skridskor.
Mannen bär en svart skjorta och hatt och ler.
En svart hund med röd krage vadar genom vattnet.
Indiska kvinnor sorterar kläder.
Tre barn leker och har roligt i ett fattigdomsområde.
Fyra tjejer i en byggnad som leker med varandra
En kvinna klädd i blått med blå väskor står utanför ett fönster.
En pojke och hans bror leker med pinnar och svärd.
En kvinna med svart handväska och röd rock sitter på en betongpelare.
En person smutsar ner sig längs en lerig stig.
En man kastar en boll på en hög av block med uppstoppade djur i bakgrunden.
En pojke går över en repstruktur på en lekplats.
En grå hund som jagar en brun hund i grunt vatten.
En man skakar hand med en skyltdocka.
Äldre män som röker när de går förbi en målning av en gammal man.
En man i svart jacka arbetar på ett tak.
Tre glashissar med folk inuti.
En massa pojkar som kör bil.
Ett barn hoppar från ett inomhus klättergym, medan andra barn klättrar över andra delar av strukturen.
Den vita och bruna hunden skakar sina öron.
En liten flicka som klättrar uppför trapporna på lekplatsutrustningen.
Grupp av människor som tittar på bärbara monitorer.
Två honor, en bär ryggsäck, står över en vattenförekomst.
Person som observerar en flod med en bro som går över den.
En kvinna med svart rock och solglasögon står framför en man som går iväg med en ryggsäck.
En kvinna sitter på en stock nära vattnet.
En man i vit skjorta och Khaki byxor med en hatt på att klättra ett berg.
Ett släde-hund team arbetar hårt på denna snöiga spår.
En man med glasögon som sitter vid ett bord med en kaffekopp och flera andra föremål på bordet.
Tre män spelar gitarr på scenen.
Två barn springer längs en strandpromenad som korsar en vattensamling.
En skallig kille med svart t-shirt spelar gitarr.
Två män sparkar en gul och svart boll över ett nät.
Unga spanska flicka hoppar från betong gård delare på trottoaren.
En nödutgångskarta hänger ovanför en dörröppning där en kvinna sträcker sig efter något.
En man inspekterar noggrant takpannorna.
En man i köket som försöker ta bort lite kött han har lagat från pappersplåten.
Ett par står och tittar på havet.
En person har sina händer i en hunds mun.
Pojke hoppar i öknen medan andra tittar och fotograferar.
En man med långt lockigt hår somnade under en biltur.
En ung pojke står och stirrar på en TV-skärm.
En liten flicka pressar en liten pojke som sitter på en gunga.
Ett barn som leker i en massa blommor.
Tre män spelar saxofoner medan en man spelar trumma i ett hörn
En brun hund och svart och vit hund springer längs det gröna gräset.
Den sida av en byggnad bredvid en kyrka är målad med en färgstark Coca-Cola skylt.
En far och son som sover i sina filtar.
En kvinna som bär grått talar in i en mikrofon vid en händelse medan två män lyssnar.
Flera personer flyttar en struktur.
Ett litet barn på ett däck svingar på ett skogsområde.
Män och kvinnor som sitter bakom ett långt bord medan de pratar och arbetar på sina bärbara datorer.
En man som är inlindad i en grå wrap lägger sig ner på marken.
En gentleman driver en maskin medan han arbetar i en fabrik.
Flera damer sitter tillsammans runt ett bord.
Kvinnan får en julklapp av en julstrumpa.
En kvinna i rosa sitter och njuter av objektet hon håller.
En hona öppnar en present.
En man som försöker hålla sig på knäna.
Två hundar är vända mot varandra på ett gräsfält.
Den bruna hunden ser en svart hund ligga i det torra gräset.
En liten basebollspelare, klädd i en vit #19 tröja, träffar framgångsrikt bollen.
En kvinna tittar på en broschyr som pratar med någon, medan en kille tar bilder i bakgrunden.
En kvinna försöker sticka armvärmare.
Två tjejer förbereder sitt hem för en stor fest.
En kvinna i en grön blommad klänning håller i en behållare med garndjur.
En ung kvinna håller upp en röd och vit klänning medan två andra kvinnor ler och tittar.
Den vita hunden hoppar över en snötäckt stock.
En människa står i ett gräsfält utrustat med en typ av trädgårdsredskap som hon använder på gräset.
En man i hatt som rider på en häst.
Den bruna hunden leker i den vita snön.
Mannen i vit kostym kastar första tonhöjden på basebollmatchen.
En man i vit skjorta gör ett tal till en mikrofon.
En kvinna som uppträder på en konsert.
En grupp unga män spelar ett spel på stranden.
En man i svart utstyrsel står framför eiffeltornet.
En man i en båt i en blå skjorta och hatt har en fiskespö som är böjd halvvägs.
Fyra rockare poserar på en stubbe.
Två killar, en bär på en väska, och en flicka går nerför gatan.
En skulptör ställer sig framför sitt verk.
En man tittar på kameran när han står utanför en tunnelbaneingång, medan en flicka bakom honom pratar på sin mobiltelefon.
En grupp människor utanför en kyrka på ett bröllop.
En grupp sittande män dricker kaffe runt två bord.
En stor grupp människor på en fest.
En man som bär brunt är ute bredvid en cykel
Folk utanför ett hus i snö.
En person som sitter bredvid ett stativ tittar på båtar i en hamn.
En man jonglerar på stranden.
En fluffig vit hund som springer över snön.
Flera personer möttes i en session, en del med datorer, en del behövde stå.
En man på en båt docka tittar på vattnet vid en båt
En kvinna i rött är något böjd bredvid en tegelbyggnad.
En man med tatueringar ligger på en soffa och håller i en penna.
Två husky-liknande vita hundar är ute på snö.
Ett barn i blå sovoverall leker med en röd mopp i en röd hink.
En vit hund som springer i snön.
Fotot tittar ner på en gata där fem fotgängare går.
Flera personer med bagage, förlorade blickar på sina ansikten, och bekväma.
Många män och kvinnor njuter av ett utomhusområde.
Två pojkar tittar på en tredje pojke som sparkar lite snö.
En man i långärmad brist skjorta sitter på en orgel i en stor byggnad som människor 3 människor ser på.
En man spelar provisoriska trummor på vita hinkar i snön.
En pojke med en tröja med dragkedja spelar franskt horn.
En man sitter med sin musikställning framför sig.
En brun och svart ner med en blå krage nära en fotbollsboll på ett gräsfält.
En man på en cykel rider förbi en klarblå dörr.
En stamman gör sin väg upp ett träd med sina fötter och händer.
En grupp mödrar sitter och ammar sina barn.
Två kor står framför folk som åker buss.
En man sitter på en bänk på en tunnelbanestation.
En man med en grön jacka och en svart hatt som står nära en dörröppning.
Den grå och vita hunden går på grus.
En man på en skateboard hoppar i luften med den.
Två manliga fotbollsspelare vilar för att ta en drink.
Ett litet barn som går genom en gammal byggnad i en blå outfit.
En hund springer genom snön.
Ett barn i blå jacka och hjälm sitter på en skateboard.
Två män jobbar på att bygga ett hus.
Barnet står på toppen av en snöbank med armarna utsträckta.
Två unga flickor i snygga klänningar står utanför.
En leksak lego finns i förgrunden medan en kvinna och barn leker med den i bakgrunden.
Ungar bildar ett rockband.
En grupp på sex personer slappnar av i vardagsrummet och spelar ett brädspel.
Surfare fånga en bra, djup klar blå, våg.
En man som står högst upp på en plaststols öga och tjurar på olika hattar
En man som jobbar på att lägga ett nytt tak.
En flicka i en badrock med en tallrik mat står bredvid en pojke som håller i redskap och en röd kopp.
Två personer sover på en bänk.
Två män och ett barn använder en linjal på en vägg.
Indisk man med elefant och grupp av indianbarn i templet.
En pojke har ett spikat armband och en konstig handske på sig.
En man som kallas Deleon talar på en Q&amp;A.
En man med glasögon talar i en mikrofon omgiven av en grupp människor.
Ett litet barn leker med en Batman leksaksbil
En kvinna som bär en grön tröja sätter godis på en hylla.
Två barn kramar varandra.
En stor skara människor tittar på scenen när en utomhuskonsert äger rum.
En liten flicka som tittar på ett stort stenblock
En svart hund leker med två mjuka leksaker framför en öppen spis.
Att se till att en korrekt redovisning av allt jag ser här registreras på lämpligt sätt.
En man tittar genom ett mikroskop medan en annan man i bakgrunden också tittar genom ett mikroskop.
En grupp killar som simmar i röda koffertar.
En svart hund med blå krage springer genom snön.
En kvinna tittar på konst i ett galleri medan två barn sitter på golvet.
En vit kvinna i röd klänning som hjälper en svart brud till hennes vita brudklänning.
Många människor nära en korsning i en upptagen stad.
En man i kostym pratar med en tjej i en blå luva i ett konferenscenter.
En man går på stranden vid soluppgången.
En grupp människor tar en promenad på stranden vid solnedgången.
Sju barn hoppar på en gräsbevuxen äng.
En beige hund och brun hund i snön.
En man som sover bakom en byggnad.
En man som klättrar på en isig glaciär med hjälp av en pick.
En liten flicka som åker skateboard medan en pojke gungar en leksak mot henne.
En man som bär en rutig skjorta målar på ett stort lakan.
En man skriver ner något bakom en buske.
En man rider på en enhjuling längs trottoaren.
En kvinna schamponerar och mannens huvud i en hårsalong.
En kvinna med blå hatt fotograferar i ett område täckt av pensel.
En brandman sätter träblock under en krossad blå bil.
En brun och svart hund som springer genom ett gräsfält
En vuxen hane knäböjer på taket och reparerar
En man visar en kvinna hur man använder en såg för att klippa en bräda.
Två personer går nerför en stad gata på natten
En grupp killar som jobbar på en liten blå öppen topp racing fordon.
En brandman arbetar vid en brand.
En vit hund springer genom snön.
En man som spelar ett svart flygel.
En ko ligger på en gångväg mellan två räcken när en del människor kopplar av i närheten och en kvinna går sin väg.
Folk med röda bygghattar som står runt en oljepump.
Två män i kampsportkläder knäböjer inför vapenräcken.
En brun hund leker i snön.
Det finns en byggarbetsplats med en grävsko och en man med spade.
Två män med ljusgula västar sitter i ett fordon.
Det finns två män i gula västar som arbetar i en stor grön fil.
En liten flicka cyklar.
En man med tunt skägg och brun jacka spelar "Guitar Hero" i ett trångt rum.
En ryttare på en häst som landar från ett hopp.
En man med glasögon pratar med en grupp vänner.
En dam med en rosa huva tar en video av stor skärmbild av ett sportlag.
En dam klädd i svart rock, jeanskjol, svarta stövlar och svart handväska, går förbi en stor annons av en dam som gräver sig igenom sin handväska.
En kvinnlig dansare gör ett språng över en scen.
En brun, svart och vit hund är på en hinderbana.
En skateboardåkare som gör ett trick på en ramp
Två förtjusande barn som var mycket lika sin mors kläder njuter av en tågresa.
En muskulös man i badbyxor spelar paddelboll på stranden
En lockig man pratar eller kanske diskuterar med en blondhårig man framför ett bord.
En polis sitter i en skåpbil och tittar ut genom fönstret.
Två män jobbar på ett cirkulärt fönster genom att stå på stolar.
En blond kvinna i blå kläder spelar cello.
En kvinna sitter i en stol medan en man tar av sig sitt strumpeband
Flera hundar grupperade tillsammans i en vintermiljö.
Den här unge mannen rakar sig framför en spegel.
En man som bär en blå skit står upp och pratar.
En indisk man som bär turban går längs en trottoar.
En man klättrar upp för en sten.
Flera dansare gör benlyft på scenen.
En skjortlös hane rider en skateboard och utför ett trick.
En japansk man i röd skjorta, på Olympics spela tennis.
En man kastar bowlingbollen för att slå ner den sista pinnen.
En kvinna klädd i en traditionell wrap kan ses genom ett litet hål valv.
En kvinna som bär en skål på huvudet går framför ett barn utanför.
Två kockar försöker komma på hur man lagar maten.
Flera män går och står i John A. Noble anläggning.
Ett barn leker bland en flock fåglar i parken.
En matleverantör som säljer mat på en gatumarknad.
En asiatisk kvinna i svarta kläder sitter på en offentlig plats.
Byggnaden är täckt med röd &amp; svart graffiti.
En man i en kanot paddlar medan en annan man kastar ut ett nät i en stor vattenförekomst.
En normal solig dag i en stor stad.
En stor svart hund blottar tänderna medan han springer genom snön.
En man blir attackerad av en schäfer.
En kärleksfull kvinna som knäböjer nära 3 katter samtidigt som hon tar hand om och matar en skadad katt.
En stor man spelar gitarr på scenen.
Ett litet barn sitter i en gunga på en lekplats.
En man tittar på ett objekt genom ett mikroskop.
Tre ljust rånade flickor sitter på en berggrund framför en stor sten.
En bunt barn går över snö.
Många människor väntar tålmodigt på att linjen skall gå ner för att komma in i denna byggnad.
En fiskare på ett fält nära en sjö.
Två små barn leker med en tonårsflicka som har ögonbindel.
En man som plockas upp av sina lagkamrater för att fånga bollen.
En ung pojke sparkar en fotboll med en ung flicka i bakgrunden.
Två lag slåss om segern!
En snowboardåkare tar en bild framför några träd.
En man i jeans och en långärmad huva, och en ryggsäck, går i en öken.
Tre unga kvinnor omfamnar medan de visar bakverk i köket.
En pojke och flicka springer över ett gräsfält mot en skogbevuxen kulle.
En grupp män och kvinnor samlas runt ett konferensbord.
Två mörkhåriga tjejer är i publiken.
En kvinna som bär en gul jacka åker skidor nerför en snöig kulle.
En kvinna står med en iller och en hund.
En hane sitter vid ett bord med en kaffekopp framför sin vänstra arm.
Ungar leker i en uppblåst lekplats.
En ung pojke svetsar en bit metall medan han skyddar ansiktet.
En man som går 3 dalmatier längs en solig gata.
Dessa tre män joggar åt samma håll längs en gata i solglasögon.
En grupp kvinnor tävlar i roller derby.
En broenhårig kvinna som bär en svart rock med kaffe i handen
En liten pojke plågar en tallrik.
Den stora bruna hunden paddlar i vattnet.
Två män i affärskläder som står bakom en kamera.
Unga vänner i en park koppla av och njuta av samtal med varandra.
Ett asiatiskt band i en parad med ett kvinnligt band majorette.
Tre flickor klädda lika i rutiga kjolar och hattar, gröna tröjor och blå knästrumpor går tillsammans.
En flicka som kastar en fotboll medan hon sitter ner.
En tjej i rosa jersey och gröna knä höga strumpor sparkar en fotboll.
En flicka som går framför ett fotbollsnät under en match.
En man, som bär en svart keps och en mestadels grå luva, verkar vara på en fest.
En man sitter på en svart och brun hund.
En röd cabriolet kör längs vägen och stoppas av en åskådare.
Svart man målar ett tecken.
En pojke som bär grön skjorta hoppar framför en fil i en bowlinghall.
De två kvinnorna tittar på något.
En tjej sparkar en boll med tre tjejer som gör samma sak i bakgrunden.
En liten flicka som spelar i en fotbollsmatch.
Fyra unga flickor i gröna och blå uniformer spelar fotboll tillsammans.
En ung flicka förbereder sig för att sparka en rosa fotboll.
En tjej fotbollsspelare står nära ett stängsel och kastar bollen tillbaka in i leken.
En äldre man som sitter ute i solen och tittar på något under sitt paraply.
En ung man och en äldre man sitter på en rutig kärleksstol.
Två kvinnor med barn som pratar med varandra.
En blond-hårig liten pojke ser framåt medan en blond-hårig kvinna justerar sin krage.
En kvinna klädd i svart är silhuetterad mot en moln mörk himmel.
Ett barn med älg på tröjan leker med ett tågsätt.
Ett barn ser nervöst ut på toppen av en bild.
En fotbollsmatch spelas när solen går ner.
En ung pojke som bär mr Potato Huvudtänder och glasögon.
Flera människor står på scenen med armarna upphängda i luften.
En flicka i gul jacka som sitter på ett stenlejon.
4 personer står bredvid en brand matlagning en måltid
En ung flicka som jagar en anka med bröd i händerna.
Två personer är tillsammans och en av dem använder en mikrofon.
En man med glasögon som klättrar upp på en stenvägg.
En man i en gul reflekterande väst knäböjer på en gräsmatta medan han använder en mobiltelefon.
Fem cricketspelare ligger på gräset.
En vit kvinna kastar upp en pojke i luften.
En ung man bär hatt och skyddsglasögon när han åker snowboard.
En man i en snorkel simmar i vattnet och tittar på vattenlivet.
Några afroamerikanska unga vuxna spelar volleyboll.
En man bygger ett stort sandslott på stranden.
En man på Rollerblades glider nerför en parkstig.
Två valpar leker i det gröna gräset.
En asiatisk man bär ett barn i en matchande morgonrock.
En man spelar gitarr i ett svagt upplyst rum.
En hund hoppar för att fånga en frisbee.
Två killar och en kvinna som står och pratar på en lekplats.
En ung flicka ligger i en snögrotta
En kvinna i blått sitter på en trottoarkant bredvid blå räcken framför havet.
Folk går nerför en gata.
En grupp unga pojkar i röda dräkter kommer med sina krukor för att fyllas med vatten.
En professionell simmare racing till mållinjen.
En man är i en pool och gör sig redo att börja ett lopp.
En indisk kvinna som använder en remskiva för att skaffa en kanna.
En grupp synkroniserade simmare ordnar sig i stjärnform i en pool.
En brun hund som skakar av sig vatten.
Två kvinnor på en film som granskar film
En man och en kvinna som skrattar.
Tre flickor bär halmhattar och dansar på en scen.
En man i träningsoverall läser för en kvinna.
En ung man och kvinna sitter vid ett middagsbord med mat framför sig.
Två glada människor går nerför stadens gata.
En kvinna böjer sig fram för att ta hand om sitt barn i en gul jacka.
En kvinna går och släpar på en resväska.
En man som hoppar i sanden längs stranden medan han håller något i handen.
Byggnation i staden på natten.
Två poliser i ljusa gula uniformer står och pratar med varandra.
En svart man drar i en blå skjorta medan han är distraherad.
Två män i kostym diskuterar ett ämne medan de står framför ett podi.
En dansföreställning pågår inför en publik.
En grå och vit pöl slåss bredvid en annan svart och brun hund på en säng.
Man i solglasögon och läderjacka tittar ner
En ung pojke klättrar uppför en spiraltrappa i ett rum fullt av böcker.
En ung pojke gungar ett slagträ på en stor baseball.
En man och en kvinna dricker vid ett bord.
En man sätter upp utrustning för en rockshow.
En person går sin hund på koppel medan ett barn i en röd skjorta rider förbi på en skateboard
En man lutar sig mot en byggnad nära en livlig gata.
En butik med Wii-konsoler i och folk som tittar på dem.
En svart hund fångad i mitten av jump fånga en leksak i munnen.
En kvinna i en rutig rock står framför tvättmaskiner inuti en tvättomat.
Män bakom fönster med galler på.
En man på en stor bit snö som håller i ett rep.
En kvinna öppnade glatt sin gåva och upptäcker en KitchenAid mixer.
Crowd väntar på Main Street tunnelbaneplattform för ett tåg.
En man och en kvinna väntar på sin mat på en restaurang.
En man med svart hår och glasögon håller en kamera på ett stativ.
En man med blå byxor i luften.
Två män i ett band spelar gitarr och sjunger på scen.
En tjej som klättrar på ett länkstängsel.
En medlem i ett band spelar ett tangentbord.
Bellingham High School-bandet uppträder.
Två män och en kvinna står i vattnet med en gyllene retriever.
En afroamerikansk man som håller en gitarr och tittar ut genom fönstret.
Barn i blå skjorta ler om vad han har i handen.
En person i gul skjorta sitter på en trottoar.
Det står en flicka på piren som bär en blå skjorta och håller i ett fiskespö.
En blond tjej sover på en soffa.
Den bruna hunden jagas av en svart hund medan han håller en liten leksak i munnen.
Två svarta och bruna hundar som tittar på varandra.
En skara människor sitter vid runda bord i en bankettsal.
Två kvinnor som bär öppna tåskor kör motorcykel.
En tjej som cyklar med hjälmen på med mulet väder.
En grupp människor roar sig vid ett bord.
En man som spelar gitarr medan han står framför en mikrofon och sjunger.
Den här damen sjunger på en klubb.
En svart hund är vänd mot en brun hund i ett öppet utomhus utrymme.
En kvinna i rosa går under tvillingflugor
Två personer i färgglada kläder hanterar fyrkanter av tyg med färgglada mönster.
En ung flicka i en beige klänning som springer nära ett skogsområde.
Två barn leker på sängen med fjärrkontroll.
Barn som spelar fotboll, en som är i färd med att sparka bollen.
En korthårig brunettkvinna som sjunger in i mikrofonen på scenen med sitt band.
En grupp kvinnor i matchande uniformer, varav en talar.
En man i svart skjorta sjunger in i en mikrofon.
En brandman dukar en röd lastbil som röker när en polis närmar sig.
En grupp människor som väntar under motorvägen.
Ett nygift par står framför en stor skara.
En grupp pojkar leker på en strand.
Två personer blir genomblöta av ett vattenfall.
Ett ungt nygift par skär upp sin bröllopstårta som de får ta emot.
Några människor sitter ner och ser en kvinna presentera något i ett klassrum som en gentleman ser motvillig ut i bakgrunden.
En barfota kvinna i en röd och grön kjol är omgiven av lerkrukor och arbetar med lera.
En pojke leker med en skruvmejsel.
Ett barn som bär en grå tröja håller en krabba och tittar på den.
En flautist spelar flöjt i ett marschband
Grabben kör sin gröna och svarta cykel nerför gatan.
Två män hänger på rep över ett vattenfall.
Fyra kvinnliga passagerare väntar på sitt tåg, en sitter och resten står.
Tre hundar springer sida vid sida på gräset.
En kvinna i grå skjorta och svarta Capris springer längs en väg.
En pojke simmar i vatten.
En man med långt hår och en grön randig skjorta talar till en kvinna som lyssnar uppmärksamt.
Kvinnor som poserar i ett fånigt foto i en studio
En ung flicka hoppade ur sin gula gunga.
En liten flicka i rött är nere på isen
Ett litet barn som är uppblandat och gör sig redo att gå ner i en rutschkana.
Flera hundar bär en man med hjälm genom snö.
Ungt afrikanskt amerikanskt barn med pärlor i håret som tittar på kameran och täcker hennes mun med en rock på.
En man lär tre flickor hur man spelar ett instrument.
En ung barbröstad man som pratar med en lättklädd man längs en ensam ökenväg.
Brun och vit hund som leker i gräset.
En kvinna i en blommig mönsterklänning använder en vävstol.
Två män i blå kläder sitter på en båt.
Tre arbetare håller hinkar och hukar på balkar med utsikt över en stad nedanför dem.
Hanspaniska människor sitter på stranden i sanden och pratar i telefon.
Ett barn hoppar upp nära en vattensamling.
Ett barn tittar på ett barn som sover i en spjälsäng.
Ansiktsfull man i kostym öppnar plånboken medan en yngre dam i formella kläder skrattar med honom.
Män låser upp en grind för ett tåg.
Kvinnorna ger mannen en kram och kyss medan hans hund är i koppel.
En man som får klippa sig i en frisöraffär.
En man inspekterar uniformen för en figur i ett östasiat land.
En ung pojke som klättrar.
En man klättrar med spanare nedanför.
Två små barn som håller varandra i handen när de går på en gata.
En svart hund som sköter svarta och vita valpar.
En ung kvinna som hoppar upp från golvet.
En grupp män klädda i rött spelar trummor.
En sidobild av Applebees och Daves och Busters restauranger.
Ett litet barn som ler på en gunga på en lekplats.
Medelålders man i gul skjorta stående på trottoaren håller en grön väska och kastar en skugga.
En kvinna med en blå halsduk läser en tidning framför en målning av solrosor.
En man och en kvinna som kysser utomhus.
En liten flicka som spelar gitarr, några blommor till vänster.
En kvinna och ett barn som båda bär röda kläder går upp på en gata
En man i en blå rutig skjorta går bakom folk med sin hund på stranden
En flicka inuti en lång tubulär bild.
En man står i fjärran på havet medan han står på en liten båt.
En svart och brun hund bär en röd leksak i munnen.
Ett litet barn går längs sidan en stor svart och brun hund med snö på marken.
En man i grå rock talar in i en mikrofon.
En grupp ungdomar som håller i flaskor och pekar på kameran.
Två kvinnor går nerför den trånga gatan.
Den lilla flickan i den rosa toppen springer nerför stigen.
En kvinna i svart skjorta som föreläser.
Det finns en liten flicka i en rosa hjälm som rider sin rosa cykel längs en vattenväg.
En banidrottare hoppar ett hinder.
En hund hoppar när han vänder sig om på en strand.
Ett band spelar på en liten scen.
En flicka i svart hatt med en rosa blomma på den spelar tangentbordet.
En familj förbereder middagsbordet för en fest.
Några personer sitter på en brygga och tittar på en sjö.
Ett band som heter Screaming Orphans håller på att ge en konsert.
Vi sjunger den populära sången för er alla.
Barn tävlar runt en gokartbana med vuxen övervakning.
En liten kropp i orange skjorta håller ett gult svärd och håller det mot kameran.
Unga pojkar som spelar boll på stranden.
En man sitter i en stol med foten uppstoppad på ett skåp och pratar in i en mikrofon.
En man i kostym sitter och pratar i en mikrofon.
En man i grå kostym pratar framför en mikrofon.
En man petar ut sin från ett litet fönster.
Någon leker hopscotch på ett utsprängt rutnät på marken.
Ett litet barn tittar på när en man spelar elgitarr.
En kille och en flicka tittar på en person som håller tal medan de sitter ner.
En man paddlar en båt under en solnedgång.
Fyra barn i svart och röd hatt och svarta kläder uppträder.
En kvinna som sitter i stolen diskuterar ett ämne i en mikrofon.
En man i vit skjorta och blå shorts som svingar tennisracket.
En pojke skär en volt i gräset.
Framför en asiatisk affär vilar en man i en stol medan en annan man städar.
Den unge pojken lekte med sitt tågsätt.
En man håller ett barn medan de ler mot varandra.
Folk går nerför trappan genom dimman.
En grupp indianer står bredvid ett gatuljus på dagen med moln ovanför dem alla.
En brun och svart hund som springer genom en flod
Människor bredvid en röd, vit och blå varm luft ballong som är på gräset
En man som talar direkt in i en mikrofon
En pojke som bär en blå huva håller ett litet djur och ler.
En grupp teaterelever hoppar i sekvens på scenen.
En liten baby i vinterkläder hålls upprätt för att ta en bild.
Folk i en folkmassa bakom en gul metallport.
En ung pojke sparkar en fotboll medan sex andra spelar men är klädda som domare.
En ung flicka klättrar på en trästruktur.
Tre hjälmbärande rullskridskor är bredvid en skridsko ung vuxen.
Två barn leker på en lekplats.
En kvinna som fixar sin dator medan hon visar sin dotter vad den gör.
Två kvinnor och en officer som avgår ett flygplan.
En man i röda badbyxor på en båt i vattnet.
En ung pojke som sover efter att ha lekt med sina vänner.
En liten flicka som bär en dekorerad hjälm är nedsänkt över en liten tvåhjulig cykel.
En man med ansiktsmask sitter nära ett tält och en husvagn.
En pojke klättrar på en blå vägg medan en vuxen tittar bort.
En arbetare som städar en tegelgata.
Den hejarklackstruppen för ett professionellt basketlag utför en rutin.
En man som tittar ut genom fönstret.
Människor framför vattnet, 3 personer sitter ner vända mot varandra som en ung pojke springer och 2 personer går mot vattnet.
En man i grön skjorta med hängslen som pratar i telefon medan han sitter vid ett bord.
En man i vit skit och beret bland många guldföremål.
En svart hund som springer i ett lopp.
Flickan i blå shorts sitter på en trasig stubbe.
Folk, utanför, kastar saker över dem.
En ung man i en blå huva som gör en vändning av en halvvägg som är täckt av graffiti.
En pojke hoppar över en annan pojke på en studsmatta.
En man i glasögon och en kvinna i svart hatt och mörka solglasögon sitter tillsammans på ett tunnelbanetåg.
En pojke är säkrad mellan två bungelsträngar och svävar i luften.
En gammal kvinna i lång rock med en liten vagn korsar gatan medan en annan kvinna röker en cigarett klockor.
En man sätter sig i en röd bil.
En ensam man kastade en fiskelina i vattnet vid solnedgången.
En man svetsar i en gul bil.
En flicka i svart sitter på golvet i en sovsal och gör klassarbete, och en flicka i röd skjorta arbetar på datorn.
Barnet är på en gunghäst av trä.
En kvinna med lockigt hår i svart jacka, svarta byxor och svarta klackade stövlar går nerför gatan.
En kvinna formar lera på en lerbrunn.
Två barn springer nerför en trottoar framför en byggnad.
En hund som kommer från en sjö.
En stor vit hund och en liten svart hund sitter i snön.
En blond kvinna skrattar.
En kvinna sitter i ett väntrum och läser en tidning som skildrar en lättklädd man och kvinna.
Någon sätter på en sko och lämnar i en hast.
En svart och en vit hund leker med en rep leksak i en bakgård
En livsmedelsbutiksarbetare knuffar flera korgar på en gång.
En äldre man som sitter framför vad som verkar vara en dörröppning.
En mörkhyad man knäböjer framför en tallrik mat.
En kvinna pratar på sin mobil medan ett par sitter på en restaurang.
Flickor i lila asiatiska klänningar sitter i stolar i en formell miljö.
En pojke i en simbassäng, bär glasögon, ger "två tummar upp"-skylten.
Ett barn springer barfota över en svart parkett.
Killen med långbrunt, lockigt hår och glasögon, spela gitarr, sitta på gräs, bära randig skjorta och blå jeans.
En kvinna som sitter mot en vägg bakom en glasruta.
En hund springer genom en skog på vintern
Folk tittar på två killar på motorcyklar.
En grupp människor står utanför och ser på när något händer.
En kille och en tjej som spelar brädspel på golvet.
En liten hund hoppar genom luften över ett snöigt fält.
Grabben med en papperskrona sitter i en kundvagn.
En man som hoppar över lådor för att träna mitt i en high school-bana.
Motorcyklist går in i en motorcykelbur framför en stor publik.
En liten flicka på en studsande lekplats djur sitter medan en kvinna tar sin bild.
En man sitter upphängd på en kursrock med en vit tanktopp.
Flera hundar går runt på en tegelgata.
En kock i köket lagar mat
En flicka med ryggsäck och en pojke på cykel står på en korsning.
Små barn leker i en hög med toalettpapper.
En äldre man sitter i en stol medan han tittar på en tidning.
En kille i kostym med en blå randig skjorta.
Folk sitter på pallar i en klädaffär.
Två vandrare klättrar medan en poserar för en kamera.
En brudtärna i en ärmlös svart klänning som håller en bukett med röda blommor på ett bröllop.
En gatuartist som spelar ett slagverk framför en skara människor.
Någon hoppar över stranden i ett tecken på glädje!
En grupp människor som sitter vid ett bord.
En pojke med hatt och shorts sover på en bänk.
En man går förbi en byggnad med en dörr där det står "Håll dig undan".
En person går bakom några ankor på vattnet till en sjö.
Flicka som spelar flöjt när hon går förbi stängsel på landsbygden.
Den vita hunden hoppar över en ström av vatten.
En dam med glasögon och en varm hatt ser på avstånd.
Ett barn med blont hår svänger på en däcksvinge.
Deli man skär kött tunn och väger de skivade bitarna.
Två personer som sitter under ett blommande träd och tittar på ett berg nära ett skjul.
En person rider i en båt på en sjö.
En kvinna med en tanktopp och handskar som tvättar fönstren ovanpå ett tåg.
En man i poloskjorta som läser för ett litet barn i knät.
En vit hund brottas med en svart och brun hund på det gröna gräset.
Två barn går upp för en enorm trappa.
En liten pojke i röd och vit randig skjorta och shorts sitter bland stora växter.
En pojke och en kvinna är på toppen av stora stenar vid solnedgången.
En kvinna i svart skjorta jagar en liten pojke i orange skjorta.
Ett barn i en röd jacka jagar duvor.
En kvinna gör ett ansikte som ser ut som hon har ont medan hon håller bröstet med båda händerna.
Två hundar springer runt i ett uterum.
En äldre man i en uttorkad fedora ler något för kameran.
En hund springer vid vattenbrynet.
Fyra män arbetar med byggnadsställningar, två har röda rockar.
Barn leker på gungorna i en park.
Ett barn och en vuxen, som var och en bär hattar, leker vid havet.
Kvinna med headscarf och flicka i röd kostym klänning gå genom urbana området.
En man i randig skjorta rakar sig mot en spegel, och ett litet barn tittar på honom.
En kvinna i en blå topp sitter på en buss.
En man som bär en röd skjorta sträcker sig ut efter sin hatt som föll medan han går en lina.
Cyklare rider nerför en livlig lantgata.
En man med en blå jacka står utanför en byggnad med guldgrimmade dörrar.
Ett stort skepp på vattnet i skymningen.
Ett par står bredvid ett stängsel och tittar på en vattensamling.
En man i kostym och slips sparkar ihop klackarna.
En grupp människor spelar tennis på en lertennisbana.
En man väntar på att få gå in i båset.
En jockey på en häst försöker hoppa stockar i ett fält.
En liten pojke i en röd jacka som glider i snön.
En närbild av en man i glasögon som tittar på kameran.
En flicka bredvid en blå presenning vägg bär en ryggsäck och en handväska.
En man med röda glasögon och vitt skägg står med käpp och träd i bakgrunden.
Barn spelar ett spel på ett fält.
En skjortlös fick i blå byxor är jagas av en flicka i en svart skjorta.
En orkester framför ett verk.
En kvinna tittar på maten hon förvarade i glaslådan.
En kvinna kramar en man utanför medan han gäspar.
En dam med grå jacka och jeans som sitter nära en man i lång rock.
En hane och en hona, båda klädda i sandaler, som går vid ett staket.
En kille fiskar utanför hamnen, det ser ut som han har något stort i slutet av sin linje.
En man i svart kostym pratar och ger upp med händerna.
En man i blått och en kvinna i rosa pos framför sjön.
En svart hund som simmar genom en flod.
En skjortlös man med en blå handduk på huvudet rakar skägget.
En äldre man försöker ta reda på vad en symaskin är.
Fyra personer i hatt står för att titta på en händelse, två av dem med kameror.
Fem personer sitter utanför och spelar kort med varandra.
En liten flicka med mörkt hår som står på en gräsmatta och samlar maskrosor.
Tre män i gula skjortor arbetar utanför en restaurang.
College män och kvinna sitter på ett möte i ett rum med en lärare medan en av männen står och förklarar något.
Det finns tre hundar som tävlar runt ett lerigt spår.
En man böjd över att sopa i källaren som är gjord för mycket korta människor.
En man sänks på en remskiva framför en byggnad.
Folk sitter i en restaurang med höga tak och stora fönster som dricker olika viner och umgås.
En lokal man som sitter på en pall visar vägen till en turist.
En kvinna i jacka står bredvid ett staket och spelar hästskor.
En kvinna i blått med en käpp sittande på en tunna.
En kvinna i röd skjorta och ett vitt förkläde arbetar med lera medan en ung flicka tittar.
En grupp vandrare vandrar längs grusstigen.
En grupp vänner som spelade en stapling spel innan det föll ner.
Den här kvinnan i shorts håller i en mikrofon.
En kvinna i svart jacka sitter på en strandpromenads bänk i trä.
En person som ligger på marken bredvid en ko.
En person sitter på gruset och håller en sovande hund.
En lycklig nygift kvinna, omgiven av vänner och familj, har en bukett med blommor.
Ett barn som bär lila rinner genom stänkande vatten medan en man i rött ser på.
Två män i ett rum med många sängar.
Två män ler mot kameran inne i en restaurang, en håller upp en öl.
Tre blonda kvinnor tittar i mikroskop.
En rödhårig kvinna sitter framför ett kedjestängsel och har två män på vardera sidan av henne.
Ett ungt par njuter av en snöbollsmatch.
Ett barn poserar med en rolig förbi för kameran vid vattnet.
En man i grå skjorta och khakibyxor sitter på en campingstol.
En ung kvinna som går i skuggorna framför ett inhägnat område.
En man som kör en kärra på en grusväg.
Två kvinnor i labbrockar tittar på en bild projicerad på väggen
En blond kvinna i en rosa polotröja hoppar med gula bungelsträngar.
En kvinna i senapsklänning med vit väska går nerför gatan framför en tegelbyggnad.
Byggande på insidan av ett hus.
En äldre kvinna och en ung pojke, som äter något, sitter mitt emot varandra.
De två sittande flickorna ler mot kameran.
Det finns två barn, en fotboll, en hund och en get ute på ett fält.
En hund med munkorg och blå jacka springer runt på gården.
En man kramar en ung pojke i en blå skjorta.
En pojke ger att vara i snön två tummar upp.
En furiös kvinnlig tennisspelare som ska träffa en tennisboll i luften.
Två personer går nerför några trappor.
Barnet i den gröna skjortan sitter på en maskin med hjul.
En man i hatt njuter av en öl.
Kvinnan tränar en vit hund att sicksacka genom metallstolpar.
En barfota flicka svänger högt på en gunga en våreftermiddag.
En polis går bort från en grind med en stor brun och svart hund.
En blond hund springer i gräset och håller en käpp i munnen.
En man står framför en staty.
En man i en allmän vägarbetares uniform sprutar vatten.
Reflektioner i vatten av människor på bro och barn promenader till vattnets kant
Kvinnan åker skridskor i parken.
Två kvinnor tittar på bilder på en datorskärm.
En rödhårig flicka har en söt get.
Ett barn som leker på en röd skoter.
Två barn, en pojke och en flicka, springer över jorden.
En person som simmar i en pool i röd baddräkt och blå glasögon.
Ett barn i drakdräkt på cykel.
En man klädd i brun rock och bombplanshatt bär påsar och går mot en korsning.
Två tonårstjejer bär snygga klänningar på ett evenemang.
Ett barn glider nerför en rutschkana medan ett annat barn tittar på
En man i kostym går nerför en fullsatt gata.
En man går framför ett äldre hem utan någon färg på det
Folk på väg hem från jobbet på tågstationen.
Två personer sitter på en bänk på en stad gata med en hjärtformad ballong i handen.
En man i svart rock och grå byxor går längs en lugn gata.
Två hundar brottas lekfullt i en stenig miljö.
En liten flicka i en solklänning leker i sanden.
En svart hund och en brun hund i snö.
En man med motorcykelhjälm vilar vid vattnet.
Sex kvinnor som visar sin nationalitet genom att hålla en flagga.
Flera personer bär vit mask håller en banner och skyltar.
Flera militärer som omger kvinnor som sitter på marken med flaggor.
Två svarta och vita hundar slåss i snön
En liten pojke leker med en basketboll och en leksak basketkorg.
Barn leker i vattenfontäner
En man med brun jacka och grå hatt står med slutna ögon i en folkmassa utomhus.
En ung pojke sitter på ett staket med ett fat mat på huvudet.
Två kvinnor med glasögon en skrattar och en ler.
En man som sitter på kanten av ett träd kantad promenad.
Två kvinnor tittar ut i en vacker skog från en avsats.
En flicka står i en affär bredvid andra butiker.
En cowboy som hänger på för ett kärt liv medan hästen under honom helt enkelt försöker lura honom.
Pojken vid poolen äter ett äpple.
En vandrare med ryggsäck går nära ett vattenfall.
Tre personer sätter upp stolar på stranden.
En man i en marin poloskjorta knäpper bilder på en golfbana medan en skara åskådare tittar på i bakgrunden.
En skoputsare arbetar när andra passerar förbi på en livlig trottoar.
En person rider på en häst i västerländsk stil, och hästen ger vika.
Gymnasieelever tittar på något och tar bilder.
En pojke och en man korsar en flod på en elefant.
En kvinna med svarta byxor och en grön skjorta jogging.
En motorcyklist med en Puma fanny-pak parkerad på trottoaren med kickstand av sin cykel upp.
En svart och vit hund med tungan ut går.
En man som sitter i en stol får håret sköljt och tvättat av andra män.
Ungar som spelar hopprep mitt på gatan.
En ung vit pojke klättrar genom en metallstruktur av stationära ringar utanför i ett stenlagt område med utsikt över en vattenförekomst.
Tre kvinnor i headscarf ser något ur ram.
Dansare övar danspositioner med varandra, och en del använder ett säkerhetsräcke för att få hjälp.
Pojken klättrar upp för en repstege.
Tjejen med den svarta T-shirten är ute med en stor brun hund.
Män utövar kampsport på bakgården.
Två kor står i närheten medan en hund ras förbi dem båda.
Två arbetare installerar en reklamskylt för en sportaffär.
En blond man, som bär en svart t-shirt spelar ett spel av scrabble och är omgiven av grönsaker.
En kamelunge går mot en kvinna, medan en man tar en bild.
En kvinna som sitter i en brun rock håller i en bok och böjer huvudet.
En man går tvärs över gatan medan det snöar.
Brun hund med öppen mun och öron i luftlöpning.
Den spräckliga hunden springer genom kärret.
En polis står vid hörnet av en byggnad.
En hund som jagar en leksaksanka.
Två barn tittar ivrigt medan en kvinna tar tag i dem orange vatten is.
En kvinna i en blå vandringströja tittar på en svart bagge.
En person i röd skjorta klipper gräset med en grön gräsklippare.
Ett barn leker nära en vältad korg med blöjor.
En man som bär hjälm har handen uppe i luften och skriker på ett liknande sätt folkmassan bakom sig.
En gul hund som springer nerför en sandig stig.
En brun och vit hund som springer genom vatten mot en leksak.
Street artist håller en kristallkula, medan en förvånad tittare tittar på.
Två små barn, en i randig topp, springer längs vägen omgiven av ormbunkar.
Hunden springer på smal grusväg.
Två små pojkar i blå fotboll uniformer använder en trä uppsättning steg för att tvätta händerna i en vuxen storlek badrum.
Tonårspojke som cyklar genom ett gräsfält.
En kvinna bär en vit väska med en röd stjärna som går på trottoaren.
Människan skyfflar trottoaren medan snön fortfarande faller.
En blondhårig tjej bär lila topp, gula byxor, olika färgade strumpor och skor.
Folk står på en tunnelbaneplattform och väntar på sitt tåg.
Två små pojkar kör förbi vuxna i sin leksaksjeep.
En man på scenen när folk tittar på honom och viftar med armarna.
En svart och brun hund springer genom skogen.
En röd bil har rullat över på en grusbana.
En skäggig man i vit skjorta och svarta shorts vandrar på en skogsstig.
Tre flickor står under paraplyer före en scen.
Den bruna och vita stora danskan leker med två gula hundar i gräset.
De två hundarna hoppar runt.
Brun hund, med grön och lila mantel, springer på gräs.
Tre ungdomar sitter utomhus och arbetar med elektronisk utrustning.
En ung pojke i orange skjorta ler när han springer på en stadsscen.
En man lutar sig bredvid en ko på ett gräsfält.
En hund som simmar i vattnet med en käpp i munnen
En man i affärskläder står i ett gathörn.
En brun hund hoppar över en gräsbevuxen hög nära en sjö.
Två män tittar ner på en annan man som står på en oavslutad gångväg.
Någon entusiast klättrar ett torn för en bättre look.
Familjen går i skogen.
Ett barn i en röd jacka pekar på vackra orange blommor.
En kvinna och ett barn äter (en picknick).
En livlig gata med två män med blå väskor.
En Oklahoma fotbollsspelare stående
En fotbollsspelare bär en jersey wuth numret "4" på den.
En fotbollstränare har ett headset.
En man springer på fotbollsplanen och bär bollen framför domaren.
En fotbollstränare tittar på en pjäs som görs.
Oklahoma Fororers fotbollslag diskuterar sitt spel medan fans hejar.
Två fotbollsspelare försöker tackla en spelare i det motsatta laget.
En leende dansare klädd i rött är på fotbollsplanen med fans i arenan blekare bakom henne.
En kvartsback gör sig redo att kasta fotbollen.
En fotbollsspelare från OU pratar med tränaren om spelet.
Två hejaklacksledare sitter på en fotbollsmatch.
En fotbollsspelare i en röd tröja får sitt knä tittat på av en annan man
En man i en Fororers jersey blockerar ett försök till UW-laddning.
Två fotbollsspelare försöker avancera bollen mot en skulle vara tacklare.
Fotbollsspelaren försöker springa ifrån motståndaren.
Fotbollsspelaren springer med bollen som spelare i motståndarlaget tar tag i benet
En hästmaskot ger high-fives till några fotbollsfans.
Fotbollsspelare på planen som en förföljare försöker ta itu med en spelare
En publik står och hejar på en fotbollsmatch.
En man som spelar fotboll som fans från motståndarlagets klocka i bakgrunden
Mannen i den grå skjortan har en blå keps på sig.
På en fotbollsplan finns det en spelare i en röd tröja och publiken är bakom honom.
En Oklahoma spelare tacklas spelar fotboll
Fotbollsspelare i rött försöker spela mot dem i lila, vitt och guld.
En grupp män spelar en college fotbollsmatch.
En fotbollsspelare som bär en guldhjälm håller i en fotboll.
Två fotbollslag ställde upp före vandringen.
Två fotbollsspelare gör en pjäs, medan det andra laget tittar på.
En fotbollsspelare springer med en boll, jagad av motståndarlaget.
De två spelarna, på motsatta lag, är mitt i en fotbollsmatch, medan andra tittar.
En fotbollsspelare tas itu med.
Två fotbollsspelare tar itu med en spelare i det motsatta laget.
En footballspelare tar itu med en motståndare.
En fotbollsspelare i rött och vitt håller upp båda händerna.
Tre fotbollsspelare bär röda tröjor är på planen.
Snacket från hans center väntar på Snap.
En fotbollsmatch pågår.
En fotbollsspelare som attackeras bakifrån av en annan spelare från ett annat lag framför en publik.
Fotbollsspelare tackla en annan spelare i en fotbollsmatch.
En fotbollsspelare för Forwards står framför oppsing laget väntar på nästa spel.
Fotbollsspelaren klädd i rött ser ner på fältet.
Fotbollsspelaren i rött sparkar av bollen.
Fotbollsspelaren gör sig redo att kasta bollen.
En grupp fotbollsspelare står bakom en coaching tjänsteman.
Huvudtränaren går ut på planen.
Ett fotbollslag som gör sina sträckor innan matchen börjar.
Många fotbollsspelare sitter på marken.
En man klädd i rött tar en bild av ett idrottsevenemang.
En Oklahoma Fororers fotbollsspelare som bär sin tröja nummer 28.
En man som bär en röd fotbollsuniform och grå handskar ser åt vänster.
En ung flicka med festhatt skrattar.
En kvinna i svart utstyrsel står i ett trägolvsrum och tittar ut genom ett fönster.
En grupp människor samlas runt en parad flyter.
En person som hoppar i luften medan han håller fast vid ett snöre som är fäst vid en stor ballong medan andra ser på.
En nybadad hund lindas in i en filt av en omtänksam kvinna.
En man och en kvinna som bär jackor omfamnar i en kram.
En man bär blå vinkar vid en busshållplats.
Ung flicka i vinterrock hoppar av ett stenblock i sanden på en strand
Flera människor väntar på ett tåg.
En liten vit hund hoppar över baksidan av en större hund för att jaga sin leksak.
En hund som bär en blå tröja har en gul leksak i munnen.
Tre spädbarn som bär solhatt leker vid vattenbrynet på en strand.
En flicka dansar som en man i kostym
Stor pälshund som går i sanden nära stora klippor.
Människor som går längs en stig längs en sjö.
En flicka med rosa randig skjorta går upp för ett set stentrappor.
En brunhårig dam i röd skjorta och svarta byxor som står och ser sig omkring.
Folk utanför på gården med två barn klättra stege till trädkoja.
En man och en flicka står framför en stor publik.
Yngre ser man bär svarta shorts och tank, med löparskor, ligger ner på en utomhus bänk.
En kvinna som går bredvid en lila vägg.
En ung flicka klädd i livfulla kläder, putsar rapphästen.
De anställda i en kulinarisk anläggning förbereda mat för att titta på kunder.
Två unga asiatiska flickor tittar ut i fjärran medan de står i ett urbant område.
En man och en kvinna står vända mot varandra framför en silverfärgad vägg.
En äldre herr som bär en randig poloskjorta som håller en liten unges hand.
Ett barn sover med sin filt på.
En man i en grön långärmad skjorta som spelar fiol i en tom hörsal.
Den bruna hunden springer i vattnet.
Två små barn sitter i identiska barnvagnar.
En gammal dam med hatt och leende.
En medelålders kvinna reparerar en del under motorhuven på sin bil.
Grupp av manliga och kvinnliga sångare på scenen.
Två män med röda västar och gröna hattar slätar ut våt cement
Män som bygger på en väg.
En man i orange skjorta och gul hård hatt går på en väg.
En byggnadsarbetare som sitter på en grön traktor.
En traktor med spade arm drivs av en orange väst bär förare på en byggarbetsplats.
Två små hundar leker på gräsmattan.
En blond dam i rosa skjorta sjunger framför en tegelvägg.
Tre personer lagar mat på köksbänken.
Några få människor och bilar ut på sin dagliga pendlande på en regnig dag.
En flicka sitter i en bil med solglasögon och hatt.
En man står i ett rött rum medan en annan sitter bredvid honom.
En kvinnlig Texas A&amp;M tennisspelare dribblar tennisbollen.
Två män i vita skjortor med matchande logotyper inspekterar motorn i en vintage röd cabriolet.
En man bankar på grytor och kastruller i sitt kök.
Det finns en man som går med en väska framför en svart fyrkantig panelvägg.
Ett litet barn på en blå leksak bär en orange skjorta.
Ett barn flyger in i ett mångfärgat ballong studsar hus.
En fet man klädd i bara shorts, parkering en röd motor scooter
Tre kvinnor joggar på en stig.
En liten hund hoppar förbi en bil för att nå en dams ansikte medan en annan hund tittar.
Ett spädbarn som bär blå kläder gråter med sin vänstra hand synlig.
Två señor medborgare pratar på en allmän gata.
En man som jobbar på en grej i ett övergivet lager.
Fyra män tittar upp på en annan man som gör sig redo att göra något.
En man som går framför en byggnad med graffiti på.
En ung man stannar för att undersöka bilden på sin kamera.
En grupp unga asiater sitter på trappan och äter och tittar på något som pågår framför dem.
En liten flicka i vit klänning som går
En kvinna klädd i en ljusgul klänning och älvvingar underhåller barn på en festival.
Tre män dricker kaffe vid ett konferensbord.
Det finns ett barn i en röd och gul leksaksbil.
Kvinna i orange jacka som leker med en svart hund
En kille som tar ett foto på en annan kille som står framför en trasig tv.
En fotograf med röd tröja är inne i en byggnad.
Fyra personer står i en tom byggnad med graffiti på väggarna i bakgrunden.
En man i röd jacka tar bilder av graffiti.
En man i jacka som hoppar runt en pinne på stranden.
En man i en kilt som spelar säckpipa.
En äldre man och en ung kvinna skrattar på stranden.
Två män spelar akustisk gitarr på en offentlig plats.
En man står i en damm och leker med vatten.
Två nakna pojkar vid en pool.
En liten brun hund med blå krage går längs en stig.
Folk blir trötta när de reser.
Två äldre damer sitter på en bänk när en gentleman går förbi dem bakifrån.
En liten pojke clowner med en colander på huvudet.
En pojke i grön skjorta håller en bild av Castro på gatan.
Ett barn som stod i gräset med armarna bredade sig.
En ung kvinna i korta ben och en tunn grön tröja går ut i en snöstorm.
En stor klippformation mitt i en skog.
En grupp människor står och pratar med drinkar i sina händer.
Kvinnan borrar ett hål i en sten täckt av blå rutor.
Två gamla män sitter framför en båt som heter Cyranka på en frodig, trädkantad flod.
En leende pojke som knäböjer i en skog.
Ett litet barn spelar gitarr och låtsas vara en rockstjärna.
Två kvinnor som håller snabbmatsdrycker skrattar.
En man med röd mössa pratar med en man i svart skjorta och en man i rosa skjorta med rakat huvud.
Tre flickor med stora handväskor går nerför trottoaren.
En man med huvudduk ger sig med slutna ögon medan han håller i någon sorts käpp.
Ett möte med ungdomar som sitter vid ett konferensbord.
En unge som bär en brun luva och gör en Ollie.
En ung person ligger i solen på en kulle och dricker en läsk.
En kvinna i tenniskläder springer för att slå en boll med sin tennisracket.
En ung pojke svänger en golfklubba med ett öppet fält framför sig.
En kvinna med blont hår ler och sätter på sig en vit tröja.
En naken kvinna dränker sig i en naturlig pool.
Två män bär en varm korg medan ett par och en man tittar på.
En tjej vattenskidor på en höstdag.
En orkester och kör förbereder sig för att uppträda framför en gyllene staty i en stor byggnad omgiven av pelare.
Två små barn under ett blått och gult paraply.
En person sitter med ryggen till en kolumn medan en annan sitter på närliggande trappsteg som leder ner.
Vit hund med mörka markeringar hoppar för att fånga ett objekt.
Pojken kommer nerför nöjesbanan på knäna.
Barn leker med träklossar i ett rum med utsikt över träd.
Tre svarta hundar leker i gräset.
En man i svart morgonrock som pratar med en annan man med en orange ryggsäck på gatan.
En blond tjej som bär en vit klänning grälar med en annan tjej med persika och vit klänning.
En man med glasögon sitter vid bordet och kollar sin telefon.
En grupp människor sitter på båda sidor av en röd sten struktur.
Två bruna hundar står tillsammans på stranden av en sjö.
En liten flicka spelar i sin leksak hus herrgård, visar flera sovrum, och några andra coola platser att utforska också.
Arbetare sköter om en byggnad med många fönster.
En stor brun hund sniffar en mindre hund i gruset bredvid en vattenförekomst.
En kvinna och två små pojkar poserar för en bild vid ett middagsbord.
En liten flicka med lila fuzzy hatt rider en trehjuling utanför.
En svart och vit hund klättrar nerför en kulle.
En grupp människor sitter i hopfällbara stolar nära tåg och tågspår.
En hund springer på ett fält.
En man som rör om i såsen med en träspatel i en stålbehållare på en spishäll.
Två hundar slåss om en grön uppstoppad leksak.
En man som sitter ner med sin snowboard bredvid en kvinna som står med skidor på ett snöigt berg.
En tonårsskateboard vid ett staket.
Två överviktiga svarta kvinnor som bär arbetsuniformer sitter på några trappsteg.
Nån med shorts och en t-shirt som hoppar över vita stolar.
En kvinna med en svart topp som står framför och håller i en mikrofon.
Två barn leker på en gård med husdjur.
Två män klädda i arabiska kläder stående i en hall.
En grupp svarta människor är klädda i afrikanska kläder, och de ser fram emot.
En ung man i jeans och jacka går nerför en gata.
Tre män står på scen och uppträder.
Två kvinnor och en man står på en scen med en gitarr i närheten på golvet.
En ung kvinna håller i en musikspelare med hörlurar när hon går.
Två män spelar gitarr i ett tomt rum.
Ett litet band som uppträder för folk på en nattklubb.
Ett fyramannaband som spelar på scen inför en del människor.
Barnen festar medan de lyssnar på sina iPods.
Fyra personer som bär förkläden och håller i en mugg i varje hand häller något i varandras muggar.
En svagt klädd kvinna dansar runt en sittande man.
En tjej och en kille som sitter på marken medan flickan blåser bubblor.
En man på en stege som skrapar lite gjutning på en byggnad.
En flicka har huvudet i ett träsnitt från ett piratskepp medan folk kastar tomater.
Tre damer är tillsammans och en av dem har 2 fingrar utsatta.
Flera dansare med tajta svarta byxor, kjolar och färgglada halsdukar dansar.
En hund springer och fångar en boll
Flera människor dansar tillsammans i synk.
En grupp sångare som provspelar på Broadwayscenen.
En sångare sjunger på kvällen på en nattklubb.
En grupp människor uppträder på scenen.
En grupp människor med vita skjortor och svarta byxor som dansar på en scen.
Folk provspelar på en scendans.
En rad flickor klädda i svart sitter på en scen.
En vit hund springer på sand.
En tjej på skidor i snö.
Man läser en tidning på en utomhusrestaurang.
Människor i en folkskara som tycks lyssna till någon som talar och kanske tillber.
En mountainbikecyklist rider i skogen.
Den lilla flickan leker med skorna av sig.
En hund jagar två gäss.
En brun hund springer genom vattnet på en strand.
En ung pojke spelar på en karusell.
Två unga pojkar som bär shorts och sandaler kastar småsten från en grusväg i en vattenförekomst.
Två kvinnor är i ett badrum och en har en kvast.
En asiatisk kvinna som ser nedstigande ut i en svart dräkt som står i bagageområdet på flygplatsen.
Barnet sitter på gräset i en park.
Här är en bild av en man med långt hår i en hästsvans som arbetar i denna statliga park.
Ung pojke hoppar från en studsmatta ner i en sjö.
Två hundar hämtar pinnar i snön bredvid trädgränsen.
En liten svart tjej som bär en blå bandanna med små guldörhängen.
En man står på toppen av ett berg och har handen på ett monument.
Två unga pojkar spelar volleyboll.
En man i kostym står på ett podi framför en publik.
En viktig äldre man håller tal för reportrar.
En kvinna i en vit tank topp sitter vid ett bord med Margarita glasögon.
En tjej i en grå skit kastar upp händerna.
En kvinna äter en måltid utomhus och sitter på en picknickbänk.
En mamma håller sitt barn i knät på en restaurang.
En man i orange skjorta funderar över sin dryck.
En man och en bebis som sitter på en filt på gräsmattan.
En man med skägg och glasögon sitter och håller ett litet barn.
En man äter en våffla bredvid ett barn
En svettig korthårig kvinna står framför en mikrofon.
En kvinna med ryggsäck sitter på en stor klippa och tittar ner över bergen.
En mustachioed man sitter som två pojkar står på vardera sidan av honom vid ingången till en gränd.
En liten flicka med rosa skjorta hoppar av en gunga.
Två små pojkar bär röda shorts och gula ärmlösa skjortor.
Två barn leker på en hög en sten.
Två fotbollsspelare båda sträcker sig för att sparka en boll i en stadion full av människor medan andra tittar i förväntan.
Man i jeans sopar den smutsiga trottoaren.
En maskerad man i blå skjorta och en slips med papper framför sig.
En man med en kamera på en kran.
Ett gäng ungar som klättrar glidande och leker på en riktigt cool lekplats.
En ung flicka utför en enhands hjul nära en liten trädgård.
Den här mannen tränar kickboxning, där det finns åtminstone en annan kille som tränar också.
En man i en lyftskopa klipper trädgrenar.
En man med orange t-shirt och hård hatt arbetar med trä-chipping maskin.
8 personer står vid en flod och hoppar för kameran.
En mörkhyad kvinna i en jeansjacka skriver något.
En man som hoppade över en vagn på Walmart.
En svart och vit hund hoppar för att fånga en frisbee på ett fält.
Två fotbollsspelare jagar efter bollen; en försöker behålla kontrollen medan de andra försöker ta den.
En kille och en tjej som pratar på cementtrappor utanför buskarna.
En nyfiken liten pojke som tittar på en snigel.
Ett litet barn som leker utomhus i en trädgård med rock och hatt på.
En kvinna visar sin ande genom att bära en lagjacka.
En svart gentleman i kostym sjunger innan en stå upp Mike
Två personer åker tillsammans på en svart motorcykel.
En man som bär grå skjorta hoppar genom luften med berg i bakgrunden.
Två svarta och bruna hundar springer genom ett fält.
Fem personer sitter i någon form av kollektivtrafik, troligen ett tåg.
Mustad man i blå flanellskjorta och brun Baltimore Ravins hatt ler.
En skateboardåkare som bär en röd rutig skjorta gör ett trick från en betongramp.
En man med en mustasch grillar hamburgare utanför.
En pojke i hjälm rider sin trehjuling nerför en gräsbevuxen grusväg bredvid ett staket.
Fyra små barn som spelar fotboll i en park.
Två små barn klädda i röda fotboll uniformer njuter av spelet.
Små pojkar spelar fotboll utanför.
Ett litet barn i sin röda fotbollsuniform sprintar under sin fars vakande blick.
Två pojkar i röda uniformer som spelar fotboll.
En liten pojke i en röd fotbollsuniform står bredvid ett fotbollsnät.
En ung pojke med bruten arm som sover i en sjukhussäng.
En grupp människor samlas för en bild medan en kvinna står på en stolpe och tar bilden.
En student använder gammal hyvel för att arbeta trä i en butik.
Två män som jobbar med en maskin i en träaffär.
En hantverkare sågar en planka av trä.
En man i blå byxor och en blå tröja gör ett räcke av trä.
En man i blå jeans och tröja fungerar
En äldre person målar en imitation av en målning som sitter på väggen.
En brun hund som jagar en gul leksak.
En man i röd jacka cyklar nerför vägen.
En man med öronskydd som arbetar på trä.
En man med orangea öronmuffar skär ett träblock med motorsåg.
En man arbetar med att bygga trappan i en byggnad.
En man spelar akustisk gitarr på en rutig säng där tre andra sitter.
En affär har bokförsäljning.
En kvinna kör sin bil med två hundar i baksätet.
En ung pojke leker på gården.
Två kvinnor som sitter ner på en fest och dricker stora glas öl.
Vissa människor ler mot varandra över några öl.
En ung man i gul skjorta och baseballhelemt som svingar ett slagträ
Man skär i en bit kött med gaffel och kniv.
En kvinna använder en linjal vid ett skrivbord för att markera ett pappersark.
En hund som väver genom en hinderbana.
Män står och pratar med varandra i ett rum med tygtak och fällbara stolar.
En grupp män som dansar utanför.
En skara lättklädda människor på en utomhusfestival
En grupp barn i fotbollsuniform jagar en fotbollsboll på en gräsbevuxen åker.
En hund som står upp på två ben med något i munnen.
En kvinna med kort mörkt hår håller i ett glas.
En kille håller en röd och vit ballong på en inomhusfest.
Fyra hundar hoppar över ett hinder.
Den vita hunden löper genom vita inlägg på en hinderbana.
En brun hund med röd krage som dyker i snö.
Ett musikbands sångare och gitarrist spelar mitt i en imponerande ljusshow.
Ett band spelar instrument för en liten publik.
En massa människor står eller sitter i en snödal.
En svart och vit hund som hoppar i gräset efter en frisbee.
En liten stråkorkester spelar i en kyrka där en publik tittar på.
Två män spelar varsin fiol.
En man utan korta och röda byxor ligger ner på en trottoar.
En ung dam som ligger på marken nära vattnet slappnar av medan hon läser en bok.
Två unga män och två unga kvinnor väntar på en buss på en japansk gata
En dam är på golvet och packar en resväska.
Människor och flera hundar i en pool i en park som miljö.
En hund, nos till marken, går på ett gräsfält.
En manlig gatuartist jonglerar en mässingsring med två pinnar, medan ett par och en manlig förbipasserande, titta på.
En kvinna klädd som en ängel sprider pappersreklam.
Folk klädda som änglar som springer nerför en gata.
En kvinna ger något till en gatuartist klädd i en vit klänning.
En man, klädd som en ängel, håller i en annan person som också är klädd som en ängel och överlämnar ett pappersark till en förbipasserande.
Två män i ängladräkter som hoppar bredvid en kvinna på kryckor.
En ung kvinna klädd i vitt med änglavingar balanserar en bowlingstift, medan en man med clownnäsa fångar en bowlingpenna.
Kvinnan bär blå jacka och orange scarf håller upp litteratur för publiken av åskådare.
En liten flicka som bär randig skjorta äter en glasskon med strössel på.
Två bruna hundar biter varandra.
En bebis kikar över toppen av en blå spelpjäs.
En man i blå skjorta står med händerna på höfterna.
På stranden stjäl en barfota kvinna i svart kjol den röda bollen från en man i gröna shorts.
En man i vit kostym som går på styltor.
Fem personer klädda mest i vitt hoppar på trottoaren i staden.
En kvinna klädd som en ängel som leker med barn.
På ett köpcentrum roar tre kvinnor i vita ängladräkter en liten flicka i svart dräkt.
Flera personer med namnmärken sitter i blå teater-stil.
Tre vuxna sitter framför ett klassrum medan en kvinna står bakom ett skrivbord.
En man i sportrock pratar in i en mikrofon.
Någon form av råd sitter vid ett bord och tittar uppmärksamt på publiken.
Flicka kysser fjäril som vilar i hennes hand.
Vissa människor sitter i en vattnig pool bredvid floden.
En man med hatt som knäböjer och tar en bild.
Damen i akvaskjorta och blå jeans sitter på en vit bänk.
Tre män vadar in i havets strand.
En grupp män som bär liknande klädryggsäckar genom landsbygden.
En långhårig man som surfar på en stor våg.
Tre män, en i blå skjorta, en i randig skjorta och en i vit skjorta pratar.
En ung man spelar flygel medan andra besöker närliggande platser.
En flicka flyger genom luften när en man står med armarna utsträckta.
En liten flicka hoppar av på en barriär.
En rocker med en blommig skjorta och slips håller en trumpinne bredvid en tröja utan trummis.
En man med pinne i fält med två hundar.
Det finns en äldre vithårig dam och en bulldog som sitter på en stubbe.
En brun hund med tunga som sticker ut och hoppar över en stock.
En tjej som åker på en cirkus som snurrar runt i cirklar uppe i luften.
En man i glasögon ber tillsammans med två andra män.
Två guldhundar tuggar en vit kudde på en uteplats i trä.
Två hundar slåss om ett tygstycke.
En person klädd i svart och röd skyddsutrustning kör en ATV på ett spår.
Ett litet barn i blå jeans glider nerför en blå rutschkana
Tre kvinnor, två med tatueringar, går nerför gatan
Hunden springer i parken.
Ett lag baseballspelare i blå uniformer som går tillsammans på fältet.
En person i rullstol är på en trottoar.
Två män pratar med en annan kille i en grön keps när en annan man sover på en bänk i ryggen.
En man i bruna kläder svänger på en golfboll med en klubba.
Ett barn glider nerför en rutschbana och ner i vattnet.
En grupp människor som går arm och arm över det gröna gräset.
En man kastar ut frisbies i luften och gränsen collie fångar dem i luften.
En äldre man spelar fiol i en bar.
En kvinna spelar gitarr framför ett träd.
Man och hopphund utföra Frisbee agera för publiken på utomhusevenemang.
En man klädd i blått som drar på ett rep som är fäst vid en båt.
En man hukar sig ner och håller fast vid sin stora bruna hund.
En man i svart skjorta och jeans står vid en mikrofon med gitarr.
En manlig gymnast svänger på ringarna.
En liten pojke med benet täckt av målare tejp, hans bror bär en superman cape.
En hund hoppar från en veranda i trä.
En ryttare på en vit häst är mitt i ett hopp över ett hinder.
En svart hund och en vit hund som leker på gatan.
Damen sätter färgat läppstift på läpparna i spegeln.
Mannen med röd skjorta hoppar upp i luften.
Två personer färdas nerför en stig som går genom en skog med ett gigantiskt vattenfall.
Overhead syn på säljare som säljer kläder och kläder.
En kvinna gör pappersmache-sfärer medan hennes vän ger sig av!
Män klädda i traditionella tyska kläder som höjer ölglas.
En vit hund följer en svart hund genom gräsområdet.
Två flickor springer genom poolen medan vatten sprutar över dem
Flickan i den ljusa röda dräkten hoppar över stigen.
En man tittar igenom produkter på en bondmarknad.
En kvinna i rosa halsduk, lila tröja, grön skjorta, håller två pojkar, båda i randiga skjortor, går i en stads park.
Två kvinnor står utanför med en ung flicka.
En kvinna håller upp en fisk som är kopplad till hennes fiskespö.
Cykling team står runt i soligt tropiskt område
En asiatisk man uppträder på en scen dekorerad med många ljus.
En kille som slappnar av i en solstol i sina solglasögon.
En liten pojke svänger i en gunga, med ett stort leende i ansiktet.
Unga flickor står på ena foten på en sten medan hennes hår blåser i vinden.
En tjej i sportkläder balanserar en fotboll på huvudet.
En kille som fyller sitt ansikte på ett möte.
En kvinna jonglerar på en offentlig plats medan hon bär en ängeldräkt.
En man ler mot en gatuartist klädd som en ängel.
Ett barn sitter i ett bad, leker med en gul leksak och en leksak dinosaurie.
En person i en blå jacka sveper upp på våt tegelsten.
En liten flicka med ett band i håret petar näsan.
Flickorna, klädda i vitt, jonglera batonger på en gårdsplan.
En gammal man med blont hår i blå skjorta och brun hatt spelar dragspel.
En hund som försöker hoppa över ett stängsel med något i munnen.
En man med en galning stående på en stege som håller gult måttband.
Folk arbetar tillsammans för att säkra en takpanel.
En man på en båt använder en stor pinne för att skjuta bort en annan båt.
En person som klättrar på en stor klippa med en annan person på marken hjälper
Ett band spelar framför en publik på en Euro Jazz konsert.
En svart och brun hund som står på en bjälke ovanför vattnet.
En man med skägg står framför en begagnad däckfirma.
Tre unga afrikanska barn i en fattig del av Afrika som cyklar.
En pojke i en surfskjorta svänger på en gunga.
En vuxen och tre barn utanför leker och har roligt.
En man håller i en liten flicka som bär randig hatt.
Pojkar släpar en apa på de afrikanska slätterna.
En man skallig, med glasögon, och en solbränd kostym jacka, fingrar strängarna på insidan av ett piano med sin vänstra hand.
Människan har fallit av en stor vit tjur i en lerig nål.
Mannen i blått poserar för en bild bredvid sin bil.
En man vadar i en flod.
En ung pojke som står på en sten bredvid en vattenförekomst med armarna utspridda.
En pojke som står på en fotbollsplan med en färgad boll.
En stor vit och svart hund springer mycket snabbt genom gräset.
En brun hund är på väg genom gräset.
En kvinna, i en t-shirt och en kjol, lutar sig framåt i ett försök att kasta en stor storlek svart boll.
En kvinna med tjockt lockigt blont hår sitter utomhus vid ett bord.
Arbetare som bär orange sliter sönder en cementstruktur med sina massiva fordon.
En man och två pojkar hoppar på en studsmatta.
En man med skägg i kaptensdräkt med cykel nästa gång.
En gul hund som hoppar från en veranda.
Tre personer står i en grupp i en park och en man läser i en park.
En grupp människor på en båt.
De tre pojkar som bär flytvästar tittar upp i vattnet.
Ett barn försöker bestiga en stor sten.
En pojke basebollspelare i en grön och gul jersey hoppar för bollen.
En flicka tränar sin vita hund med godis.
En afroamerikansk flicka som just hade fått en docka från en familj som adopterade henne från staterna.
Fyra små barn visas i denna bild med byxor och skjortor medan de sitter i rummet.
En person som vandrar uppför en kulle i snön med en hund.
En pojke hoppar ner i vattnet i den blå poolen.
Fem pojkar sitter på en grå flotte i sjön.
En man som jobbar på en byggnad tre våningar upp.
En man i en blå väst sitter uppfälld utanför ett fönster med en färgburk.
Mannen i ryggsäcken tittar åt vänster.
Tjejen springer genom ett fält med en brun hund och en vit hund.
En man och en kvinna handlar tillsammans i en stad.
En liten pojke knäböjer och förbereder sig för att kasta en basketboll.
Folk står framför en skylt där det står "Den djupa änden".
En ung kanna, klädd i en maroonskjorta och hatt, har just kastat ett kast.
En man som bär kamouflage är nere på alla fyra.
En Chelsea fotbollsspelare (Frank Lampard) och en Liverpool fotbollsspelare båda göra ett försök på bollen medan domaren tittar i bakgrunden.
En kille med glasögon jobbar på en dator på sitt kontor.
En man i röd skjorta som försöker hoppa för att få ett handtag i ett bergigt hörn.
Fyra män som drar en kanon på en vagn.
En kvinna kastar ett föremål på ett mål och försöker vinna ett pris på en karneval.
Två hundar leker i sanden.
Två män står på en brygga och tittar och pekar på båtar.
En man med orangea stövlar står med några andra människor.
En vandrande vakt står framför en asiatisk byggnad.
Njuter av en parad på en varm sommardag.
Person som står i vattnet med en gul båt med en åra i handen.
En ung pojke skyfflar sand till en form.
En svart hund med brun munkorg som simmar i vatten.
Två kvinnor sitter vända mot varandra medan den ena tittar ut genom fönstret och den andra läser en bok.
Bluffig bild av en ung pojke som knuffas i en vagn av en annan.
En svart och en brun hund.
Ett litet barn som rider på sin pappas axlar
Två kvinnor undersöker en glaslåda.
Två fotbollsspelare jagar bollen.
Sex barn springer genom ett blomsterfält omgivet av träd.
En man målar ord på framsidan av ett säljstånd.
Två barn klättrar på kedjor mellan två trästolpar.
En äldre person som bär glasögon och en överdimensionerad grå rock sitter i en dörröppning.
En kvinna i vita kläder sitter på gatan.
En man sitter nära en cykel medan folk gör val från en gatuförsäljare i bakgrunden.
En man trampar en ovanlig cykel förbi en brandbil.
En man hoppar för att fånga en frisbee, medan en man och en kvinna springer mot honom.
En grupp människor med ett tecken som säger "Maritime arbetare säger stoppa svarta dödsfall i förvar".
En svart hund och en brun hund med en käpp i munnen springer ut på fältet.
En grupp på fyra vandringar genom en snöig skog.
En kvinna och en hund med rumpan vänd mot kameran
En pojke blåser bubblor
En liten flicka blåser bubblor genom en gul båge.
Det är en man som jobbar på en skylt.
En spelare föll ner på en hård domstol i kvinnors volleyboll.
En volleybollturnering som sponsras i ett spanskt land.
En man som bär gul skjorta och bär kaffe på trottoaren
Två små pojkar håller upp skålar med mat till kameran.
Två män, en med svart skjorta och den andra med vit skjorta, sparkar varandra utan att få kontakt.
En ung flicka hoppar i sanden på stranden
En skjortlös man skrattar åt sin vän som poserar för en bild med en drink i handen.
En polis står i en dörröppning.
En solbränd greyhound som bär en guldskjorta med ett nummer på springer nerför ett spår.
En kvinna står på ett blomsterfält.
En man som spelar med en fotboll som två andra ser på i en stor utsträckning av gräs.
Rödhårig kvinna svarar på frågor när hon sitter vid ett bord för pysselzine.
En man med röd och vit skjorta och blå shorts, hoppar för att slå en tennisboll med sin racket.
Fyra personer spelar ett spel i gräset.
En man i en ugn som delar mellanmål med sina barn.
Många barn leker utomhus i gräset och övar slag.
En pojke i en blå skjorta på en hög av lera
Mat och dryck på en japansk marknad.
Ett litet barn leker med en färgglad leksak utanför.
En tjej i vit hatt hoppar för att spela tennis.
Vid någon slags stor sittande händelse gör en man och ett barn konstiga poser.
En äldre kvinna gör te i sitt kök.
Två flickor slåss på skolgården.
En liten flicka klättrar upp för en stenvägg.
En liten pojke i svart skjorta som ligger över tegelstenar och sticker handen i leran.
Ett par människor som kämpar genom en lerig grop
En man som bär baddräkt dyker ner i en pool omgiven av en skärm.
En flicka sitter på en stol i ett vitt rum.
En man sitter i en trästol framför en vit bokhylla och orange lampa.
Många motorcyklister rider längs gatan.
En person med fiskespö är bakgrundsbelyst mot en blå molnig himmel.
En man håller upp en fisk han precis fångat.
En man duckar ner mellan de röda tulpanerna på ett blomsterfält.
Ett litet barn med blå sandaler rider en skoter nära stranden.
En ung asiatisk pojke springer med en vit och grå hund på grönt gräs.
En liten pojke är i ett badrum med en grön boll.
En far och son flyger en röd drake.
En man på havet.
En ung pojke i röda Crocs och en hjälm hänger från en klättervägg.
Tre personer samlas och binder pinnar eller pensel.
En man i en keps deltar i en protest mot ICE Raids framför Stonehurst grundskola.
Vissa människor sitter runt en brand och dricker.
En ung pojke med rött hår och gråfärgade ögon sticker ut tungan.
En man som bär trä i vildmarken.
Person på en wakeboard i luften
Folk utövar kampsport i en träningssal.
Två flickor i karateuniformer kämpar i en dojo.
En man är skysurfing på vattnet.
Två lag flickor på planen gör sig redo för fotbollsmatchen.
En flicka i en röd, vit och blå fotbollsuniform som spelar fotboll.
En man i vit skjorta och klänning byxor sitter precis under en sten valv.
Personen håller en bild framför sitt ansikte.
Fyra personer sitter runt en TV och spelar ett tv-spel.
Två män stirrar på varandra och bär landsspecifika uniformer.
Två män som ser väldigt lika ut med skägg slåss om en våffla.
En man med en svart ärmlös skjorta som gör byggjobb.
En man i en mörk tank-topp håller i en järnstång medan man tittar åt höger.
En man i en svart tanktopp röker.
Medan du spelar fotboll flicka i röd randig skjorta går in i flicka i vit skjorta.
En man i röd skjorta lär sig att klättra uppför en klippa.
Buddhistisk man med glasögon sitter vid mycket dekorerat skrivbord i färgglatt kontor som viftar runt en påfågelfjäder.
En kvinna som håller en liten boll och jagar en liten pojke.
En blond hund springer nerför en stig bredvid en rhododendron.
Mannen somnade under arbetet eller klassen.
Tre personer simmar i vattnet och en person på sanden springer ner i vattnet.
En hindi man sitter bakom ett bord med en klocka tittar på objekt.
Blond flicka ler medan hon sitter på vägkanten.
En man sitter vid en brygga och tittar på vattnet.
En flicka sitter på en stenvägg medan hon tittar på sin mobiltelefon.
En liten pojke som sparkar rosa fotboll på en basketplan.
En kvinna med halsduk står nära vattnet och tittar ner.
En kraftig man på plaströren som böjer sig i en svart och vit polotröja.
En person flyger med en gul fallskärm ovanför en grön byggnad.
Barn som leker med trasig kontorsutrustning.
Tre män häller cement från en cementbil.
Byggarbetare i orange som arbetar vid en gata.
Det finns en man i en lätt skjorta som klättrar på en klippa.
En vithårig man stirrar på en metallstav.
En man ligger under en stor mossig klippa i skogen.
En svart hund stänker i vattnet.
En byggnadsarbetare i en vit hård hatt med en stamtatuering på höger arm som arbetar i en böjd överposition.
Närbild av lilla flicka dans
En brun hund som springer genom en damm.
Damen i en blå skjorta som verkar glad över tidningen hon håller i.
En grupp kvinnor skrattar medan kvinnorna med blå topp håller i en grönbok.
En sångare som sjunger för folk att höra.
De sex barnen är i skuggan av ett lummigt grönt träd.
En gul hund går längs en bergsstig
En liten pojke tittar på en Ferris Wheel i rörelse.
En ung, barfota flicka i röda solglasögon spelar i ett handfat.
Två barn delar ett utrymme som gör det möjligt för dem båda att maximera sina individuella ambitioner.
En stenskulptör som arbetar på en sten.
En man klättrar i berg vid solnedgången.
Ett barn i svart hatt och blå skjorta står bakom en trästolpe.
Det lilla barnet står i en kampsport pose.
Två båtar manövreras nerför en lugn flod.
Två personer i en båt paddlar sig förbi stora träd.
En skalle med roddare på en sjö.
Två svarta hundar leker i vågorna på stranden.
En person som hoppar i ett sten- och trädfyllt område.
En tonårspojke springer genom jorden nära ett hus på landet.
Folk samlades på en medevil-festival.
Två unga pojkar i swetashirts på en lekplats
Två personer sitter på en stubbe bredvid en bäck.
Kvinnor i vita klänningar åtföljs av män i smoking när de går in i en kyrka.
De här människorna slappnar av i det höga gräset.
Liten pojke sträcker sig efter blå bar i lekområdet, ett annat barn i bakgrunden.
Två hippies spelar musik i quad, en har till och med blått hår.
En man som rör sig ur ett hjulfat.
En man som håller i en grön bowlingboll står vid bollåterlämningsmaskinen i en bowlinghall.
Två barn som rider trehjulingar passerar en rosa banderoll.
En kvinna i rött sitter på kanten av en brant klippa.
En grupp människor både vuxna och barn står runt ett gäng får.
En man som joggar i ett maraton
Två killar som knäböjer på marken och gör en gest mot himlen.
Ett band spelar i en bar inställning
Fyra cowboys som sitter vid ett bord och dricker Jack Daniels mitt på en rodeoarena.
En liten flicka i randig skjorta ler på en restaurang.
Mannen bär svart skjorta böjd över med hjälp av en såg för att skära igenom sten.
En ung pojke och en ung flicka läser en bok tillsammans.
En kvinna väver med en kam i handen.
En målare på en stege målar tegelstenens yttre blå.
Den blonda kvinnan hukar sig på ett fält av rosa tulpaner, nära ett gräsfält och träd.
Tre magra, numrerade, gråhundar tävlar längs en bana.
En man rider en go-cart på go-cart banan.
En liten godisförsäljare säljer under ett tält på natten.
En man utför en fysisk bedrift när människor går förbi och ser hans prestation.
En grupp tjejer som sitter tillsammans och pratar.
Fyra unga barn har en bild tagen av dem i luften.
2 flickor som tvättar ett golv täckt av tvål.
Pojke i röd skjorta som står på ett plastföremål och håller i en gul leksaksskyffel.
Ett litet barn jagar vatten sprutar i en fontän.
En man med vit skjorta, svarta byxor och vita strumpor på hotellrummet har hoppat upp i luften för att landa på sängen.
En man sover på en fåtölj på en trottoar.
Flygvärdinnan klädd i gult visar användning av flytväst.
Två unga flickor som håller varandra i handen och går nerför en stig vid skymningen.
En publik tittar på en baseball match som en man gör det till basen medan en annan man försöker få bollen.
En stor hund springer på gräset.
En hane i en keps sitter på en vägg målad svart och gul.
Tre svarta flickor med vita skjortor leende
Ett barn i jacka sitter i gräset.
Flera män står tillsammans bakom ett räcke.
En äldre, flintskallig man sitter vid datorn med en reflekterande orange väst på i en arbetsmiljö.
En man på en motorcykel går runt hörnet.
En man med blå väst och bruna byxor som vandrar uppför ett berg.
Hunden försöker bita en stor blå boll.
En man i röd skjorta och en kvinna i khakiskjorta står och pratar.
En svart hund skakar vatten från kroppen.
Den lilla flickan bär en vit T-shirt med fredstecken och en havsskumgrön tutu.
En man i Seattle har en skylt som ber om pengar.
Två vänner går nerför gatan och för ett livligt samtal.
Tre män arbetar på ett hemförbättringsprojekt.
En kvinna som går till jobbet framför en familj på semester.
En hund som springer på stranden
En man i jeans och en röd rutig skjorta står inne i en telefonkiosk.
En grupp människor på en trottoar och en kvinna med städredskap.
Två män sitter på trottoaren med kundvagnar fyllda med sina tillhörigheter.
En medelstor brun hund som hoppar
Ett par händer inblandade i en uppgift.
En grupp människor i en modern och avslappnad restaurang.
Från denna vinkel kan du se kakelgolvet mönster i denna restaurang mycket bra.
Ett barn springer på en krittäckt trottoar.
Två vita hundar springer i gräset tillsammans.
Två barn går nerför en stig i skogen.
En man klädd i jeansjacka och svarta stövlar sover på golvet.
En kvinna som ska äta i ett vitt rum.
De två kvinnorna i mitten håller i röda burkar.
En föreläsning för en kvinnogrupp.
Två kvinnor som markerar ett papper medan de står i en skara människor.
Tre kvinnor tittar på ett objekt på en soffa.
Två män står på en pir bredvid en vattenskoter.
En spoof drag queen dansar på en bandscen.
Två kvinnliga hejaklacksledare gör ett jubel medan de lyfts upp i luften av manliga hejaklacksledare.
En man som håller i en flaska står över en grill.
En kvinna som säljer sina varor på filtar på marken med en stenmur bakom sig på en utomhusmarknad
En hund som simmar i en damm
En brun hund sniffar en vit hund som ligger på golvet.
En man på jobbet med en marinfärgad tröja som dyker.
En man på en motorcykel gör en wheelie på banan.
Två tunna hundar springer snabbt genom högt torrt gräs.
En brunhårig dam ler mot kameran framför träden.
En gammal man som städar sopor på gatan.
En man i skyddsväst sopar sopor på en utomhusplats.
En man som sitter vid ett bord i en restaurang.
En tonårsflicka med kort brunt hår stickas med stora nålar och grått garn.
En man som kastar en käpp för sin svarta och bruna hund.
Svart kille i svarta shorts studsar fotboll på huvudet på stranden nära vatten med en annan man tittar på honom.
Tre män arbetar tillsammans på ett fält.
Ett barn som bär ett rött ögonskydd sträcker sig ut för att röra vid en mycket stor bubbla.
En person går på en livlig gata medan han bär ryggsäck.
En kvinna i svart klänning och platta skor håller i huvudet medan hon väntar på att gå över gatan.
Tre barn drar ansikten på en lila bänk.
En mor leker med sina två barn på en såg.
En man som hoppar från en ramp på en skateboard i en fullsatt park.
En ung pojke bär däckgummi på en smutsig väg.
En man som gör sitt chip under mikroskopet
En grupp barn som poserar för en bild utanför en husvagn.
En brun och svart tjur springer från en liten svart hund.
En man gör tricks på en cykel på en ramp medan en publik tittar på i närheten.
Lokal säljare i staden säljer sin produkt till stadsbor.
Ett par kyssar på en livlig trottoar.
Folk går på en trottoar bredvid spårvagnsspår.
En mans och kvinnas trädgård tillsammans en solig dag.
En kvinna spetsar volleybollen medan den andra försöker blockera.
En svart hund springer på gården
En grupp människor går genom en karneval.
En man klädd i lila skjorta och röd bandanna ler mot dem som tittar på honom.
En kvinna med solglasögon och en blommig skjorta ser åt vänster.
Två personer står vid en kamel med behållare fastspända på honom.
En kvinna som ser barn leka på ett träd.
En skara människor som går på en trottoar i en stad.
En tjej med rött hår hoppar på en sanddyn.
Ett formellt klädd par, hon med munnen öppen, står bredvid varandra.
Några kvinnor som spelar volleyboll.
Det finns en stor publik framför en byggnad.
En man sitter på en bänk och läser en bok.
En grupp människor är utanför en tegelbyggnad och tar bilder.
Hundar som springer och leker i ett gräsområde.
En hund väntar på att en man ska kasta en boll i havet.
En pojke snurrar på en park lekplats.
Fyra män och en liten pojke som sitter runt en inomhusbrand.
En förälder håller tillbaka sin son från att hoppa på spåren.
Ett barn sticker huvudet ur taxin och skriker.
En man talar in i en mikrofon på ett podi.
En man verkar laga mat åt kunder på gatan.
Kvinna väver medan unga flicka sitter i närheten med färgglada vävning runt omkring dem.
En kvinna med en blå hatt på att hålla ett paraply med en stor publik bakom sig.
En gul hund springer genom gräset.
En hund ligger på ryggen nära ett barn och läser en bok.
Tre personer samlas på en konferens.
En restaurangmiljö inne i en byggnad där människor för närvarande äter.
Två män pratar med varandra.
En svart och vit hund hoppar högt för att få en grön Frisbee.
En svart hund som hoppar för att få en fotboll.
En man i en grön t-shirt på en lina som hoppar från en sten till en annan.
En ung kvinna skjuter mot ett mål.
En olycka med en grön Sudan och en grå skåpbil.
Ett barn som flyger en drake.
En liten pojke sitter bland andra i folkmassan med en nyfiken blick på sitt ansikte.
En liten brun hund i gräset försöker fånga bubblor
En vit hund med beige fläckar springer genom ett fält.
En man i svart skjorta håller handen av en liten flicka i flätor.
En ung pojke i en blå och brun skjorta leker i smutsen med en rake.
Rum av människor som använder datorer, och testa teknik.
En man som jobbar på en ljus orange maskin.
Tre barn leker i trädgården.
En ung man i svarta kläder går inomhus förbi en rad datorskärmar på.
En hund springer mot en boll för att fånga den.
En svart hund och en grå hund springer på stranden.
En kvinna i solglasögon som dricker vatten på flaska.
Två män sitter med munnen vidöppen.
Folk pratar på en utställning.
En kvinna gör en gest med händerna när hon sitter på ett café.
En man i ruffles knuffar en barnvagn genom en park.
Två unga vuxna stannar för att ta en bild med män klädda i kostymer.
En transvestit som står på en stadsgata i en polka-punkt-fickup och fisknät.
Kvinnan i klänning och hatt sitter på trappan med huvudet på händerna.
En brun hund jagar en frisbee
En man i vit skjorta och randig slips som håller tal på ett podi.
En man i kostym håller en presentation i en byggnad.
En grupp kvinnor som står framför en blå Sallie Mae-banner.
Gamla människor sitter och skrattar på en restaurang.
En kvinna som bär en krona på huvudet sticker ut från folkmassan i en park.
En blond kvinna och en man samlas utanför med folk.
En grupp hejaklacksledare som arbetar och planerar några av sina rutiner.
Tre kvinnor i neon baseball kepsar och hjärta t-shirt hejar.
Två bruna hundar leker med en blå leksak i ett grönt gräsfält.
En arbetare arbetar på glaset i en hög byggnad.
En gatuförsäljare läser en tidning medan han väntar på kunderna.
En brun hund springer genom gräset.
Ett leende barn med randig skjorta, som hålls av en kvinna med grått hår.
Pojke kryper genom en cementtunnel.
Barn i blå luva och shorts glider nerför en rutschkana.
En tjej som ler mot kameran från en repsving.
En ung pojke i vit skjorta sparkar en boll i ett mål.
Barn som bär hjälm rider hästar i en ring.
En svart och vit hund som går över en blå hundramp
Två hundar leker, en fångar en frisbee.
Människor som äter utanför en restaurang, njuter av sig själva och dricker öl och andra drycker.
Många människor är samlade runt staden gatan.
En ung kvinna skriver ett meddelande i krita på trottoaren.
En hund hoppar av en hund hoppar.
En kvinna håller i ett barn när hon skriver med en grön markör.
En ung man drar i ett rep medan han äter en smörgås, barfota.
En ung pojke som bär mössa håller i solglasögonen medan han skriver på en banderoll.
En afrikansk pojke sippar på sin sked i ett grönt rum.
En man som bär snorkel och goggles ger tummen uppåt när han och en annan person skyndar sig genom vattnet.
Två kvinnor skriver på ett lakan.
En rad människor har bildats under ett tecken medan andra människor ligger på marken.
En man talar animerat till en person i orangutansk kostym.
En mycket glad pojke skriver på ett stort papper med många namn på.
Två flickor sitter på marken och en bär en djurdräkt.
En kvinna i vit skjorta och lila pannband sitter och håller i en stolpe med vit duk.
En båt som seglar förbi den stigande solen.
En man med kamera och hund på en grushög.
En kvinna som bär en gul taxidräkt poserar på en gata.
Ett band spelar på en konsert medan publiken höjer händerna över huvudet.
En gammal man bär en svart jacka.
Två hundar springer genom en låg liggande vattensamling.
En skara människor som sitter utanför en byggnad.
En lätt överviktig ung man, med långt svart hår och en grön tröja, lutar sig tillbaka i en stol och håller en flaska mot bröstet.
Det här är en ung man som hoppar mitt i luften på en studsmatta.
En man i förkläde testar mat medan han lagar mat över en spis.
En kvinna i ett blått förkläde som lagar mat i ett kök.
En vit hund med orange band hoppar upp för att se en bänkskiva.
En man med cigg går förbi Graffitti som säger "Var är du?"
En ung man i en blå t-shirt håller upp handen mot munnen medan han sitter på en soffa.
En ung kvinna mitt i hoppningen på en studsmatta på en vacker landsbygd.
Barnet glider nerför en blå rutschbana med mamma längst upp på rutschkanan.
Sex personer forsar i en flod med dallandskap.
En asiatisk eller kinesisk man som sjunger en sång med inriktning på en asiatisk eller kinesisk kvinna.
Två små flickor går ut i solskenet.
Nödpersonal tar hand om ett offer som behöver hjälp.
Toddler i pyjamas leker med pappersklipp av bokstaven "P".
Två honor står bredvid varandra och tittar upp i taket.
En kvinna gör kaffe på ett kafé.
Pojken med den blå skjortan springer på gräset mellan träden.
En flicka på trä och en man som går ut.
En folksamling med folk som står uppradade framför en teater.
En man med dragspel går nerför gatan i ett offentligt område.
En äldre kvinna i stamklänning väver färggrant tyg.
Den svarta hunden fångar något grönt i munnen.
En stor brun hund springer genom ett gräsfält med tungan hängande.
En liten flicka håller vattenslangen för hunden att dricka från.
En hund som deltar i ett lopp medan han bär nummer 6.
Ett ungt par slappnar av mot en stenmur.
Två kvinnor på gröna stolar tittar på en bok.
En galen man gör stöten med en bil när en vän ser på och skrattar.
En skäggig man med röda shorts, en svart t-shirt och spegelformade solglasögon lutar sig i en fällbar stol.
En kvinna i gul skjorta står vid matstånd.
Tre unga flickor med solglasögon dansar och sjunger i ett familjehem.
Sting sjunger och spelar gitarr inför en publik.
En man i en gammal kostym som håller upp en protestskylt i en skara människor.
En svart hund bär en leksak på gräset.
Barnen är under en stor fontän i staden.
En man och en kvinna leker på tunnelbanan.
Ett barn hoppar av en gunga medan det är i rörelse.
En man slappnar av i ett badkar med vatten och ett ljus som lyser bakom honom.
Två män på en scen som spelar gitarr och sjunger.
En kvinna går nerför trapporna med en liten flicka på en arena.
En tonårspojke håller upp ett stort vitt pappersark vid ett evenemang, med två småbarn också på bilden.
En liten pojke går med en liten rosa flagga.
Tre ungdomar står på gatan och samtalar.
En man i luften som håller sin cykels styren
En svart och grå bronco försöker lura en cowboy på rodeon.
En grupp människor står runt på en gata.
Ljusblå bil går nerför en grusväg, som åskådare klocka.
En man äter majs på kokset medan han pratar med en kvinna.
En kvinna som bär glasögon håller i en spegel med ena handen medan hon ritar en bild med den andra.
Biker stannade på en väg.
En stor grupp tonåringar sitter inomhus i gula säten.
En liten pojke har en dekorerad kartong på huvudet.
Två män, båda i blått, står på en båt med en pistol.
En person äter nudlar.
En man ligger på marken och skrattar under en match.
En man som spelar cricket
En man och en hund på en strand.
Tre personer diskuterar processen för att inrätta ett socialt evenemang.
En man med mörkbrun skjorta klättrar uppför en stenig höjd.
En kvinna håller ett barn medan ett annat barn ser på.
En man i rosa tuggar en tandpetare på tunnelbanan.
En flicka i röd kjol med några hula hovar
Tre unga flickor och två blonda kvinnor hoppar rep på bok.
En racerbil rör sig längs vägen när två personer tittar på avstånd.
En man i en ärmlös blå skjorta och atletiska byxor slår en boxningssäck.
Den dränkta hunden simmar.
Folk som sitter utanför med ett stort träd på vänster sida.
Två kvinnor slåss i en kampsport turnering.
En tonårspojke i vit skjorta talar till en grupp tonåringar som sitter vid picknickbord framför en park.
En hund simmar genom vattnet.
Detta är ett barn, klädd i rött och blått, svänger på en gunga.
En kvinna som tittar ut genom ett fönster.
En man i vit t-shirt hoppar något på sin gula cykel.
Ett brudparty ställer upp för en gruppbild.
En grupp människor i gräset medan en person till höger sitter i ett träd.
En gammal man som skalar morötter framför en folkmassa.
En man och en kvinna spelar fiol utanför ett fönster.
En liten hund som fångar en boll i munnen på en strand.
Grill för tre på strandpromenaden med utsikt över vattnet.
En man klättrar stora stenar.
Den bruna och vita hunden fångar en frisbee i munnen.
En grupp människor picknick på en gräsbevuxen kulle nära havet.
En flicka i svart skjorta tittar åt sidan medan hon sitter på en träbänk.
En far och en son matar fåglarna en vårdag.
Det finns tre kvinnor i rosa klänningar som står upp och dricker ur vinglas.
En grupp människor i halvformell kläddans.
Flera människor går på gatan och man har en cigarett.
En man i skyddsdräkt tränar en polis schäfer.
Tre får betar på gräsfältet med en hund som går bakom dem.
Konstnär på gårdsplanen sitter teckning med människor i förgrunden.
Fem unga flickor framför ett grönt tält, fyra sittande och en stående, njuter av ett mellanmål och har ett samtal.
En ung flicka gör sig redo att slå en softball.
En båt med flera man dras till land av ett stort team av hästar.
Den unga fotbollsspelaren försöker undvika att angripas.
En grupp människor njuter av öl i parken.
En kvinna i blå denim shorts sitter på stenvägg.
En grupp män i en gul båt med sina hundar.
En man kastar en grön frisbee i en park.
Ett par unga pojkar i t-shirts gömmer sig i skogen med en som ser hemsk ut.
En liten pojke i en kilt fiskar med en pinne.
En flicka i vit klänning går mot vattnet och bort från vita stövlar på en strand.
Ett par kyssar i en skuggig gångväg.
Amerikansk hatt är med blå stjärnor och röda ränder, ser vacker ut på den här tjejen.
En man börjar sin dag i Indien.
Den svarta och vita racerbilen avrundar svängen.
Sex tävlande i ett mycket nära cykellopp alla i olika färger uniformer.
En brun och vit hund som leker med svart hund.
En man står i ett nedslitet område.
En man målar en gul linje på gatan.
Det finns en lockig brunett som läser en meny.
En man klädd som polis, har en falsk gam upphängd på armen.
Två gula hundar leker med varandra.
En pojke står i poolen på botten av en blå vattenrutschbana.
En vit bil racing i smuts och vatten
En röd rallybil tar en hal sväng i ett lopp.
En gul racerbil glider genom ett hörn som åskådare klocka.
3 personer, en man som spelar gitarr medan han sitter på golvet och två personer spelar ett spel på en soffa.
En ung man hoppar på ett bord.
Två basketspelare i high school sträcker sig efter bollen och en faller ner på golvet.
En man i röd skjorta med ryggsäck som går förbi en automat.
En man i grå kostym pratar med en annan man i svart kostym.
En man som sitter i en båt flyter nära en grotta.
En man i gröna skjortor sitter och designar en fällbar fläkt medan han väntar på kunderna.
En bebis som bär en blå jacka sitter i sand.
En man som bär en grå tröja och bruna shorts skär gräs med en gräsklippare.
En man i grått är en levande staty.
Den lilla flickan sitter på en gammal bänk och gör ett ansikte
En äldre man sitter bland högar av metallskrot och verktyg.
En man står på en gräsbevuxen klippa som hänger över ett djupt blått hav.
En liten pojke skålar i en mattad hall.
En ung pojke i randig skjorta som springer nerför en sanddyn.
Två långhåriga män med skägg som spelar instrument, den ena en banjo den andra en fiol.
En grupp människor står tillsammans utanför när man fotograferar.
Lilla flickan i rosa är på väg.
En kvinna bär en halsduk över håret på avstånd bakom några blommor.
Väskdamen går igenom soporna.
En grupp människor samlar olika föremål framför ett fallet träd.
Åskådare som tittar på vit och blå racerbil som passerar förbi.
En liten unge som springer ut i havet med duvor överallt.
En racerbil gnisslar genom en sväng som åskådare klocka.
En ensam kvinna i hatt sitter ute på en bänk, under ett träd.
Ett vått barn som står i vatten.
Tre kvinnor som går nerför gatan en regnig dag.
En man tränar sin kropp att dra i en tunna.
Arbetarna städar trapporna och fasaden på en stor staty i en park.
En flicka som springer genom ojämn sand med lite förvissnat gräs.
En vit och solbränd hund springer genom det höga gröna gräset.
En flicka och en pojke studsar på stora bollar.
En flicka i vit klänning som håller rosor ger lite till en man i en grå tank topp.
Fem personer deltar i en diskussion på en scen.
Tre barn leker på en gunga en sommardag
En man i glasögon tittar på sin elektroniska apparat.
Två människor hukade sig nära marken i en mörk gränd.
Flickan med röd rock går över gräset.
En kvinna med rosa halsduk pratar i telefon framför en Pink-butik.
Ryttare i ceremoniell dräkt rider vit arabisk häst, också bär ceremoniella filtar och tofsar.
En kvinna som bär en klarröd klänning och ljusröda skor går på grå trottoar.
Killen med nummer 12 jersey kastar fotboll.
En grupp fotbollsspelare som väntar på att spelet ska starta
Sex arbetare jobbar på tågspåren.
Män i orange uniformer är i en tunnel.
Järnvägsarbetare som arbetar på spåren nattetid
Hårt arbetande arbetare som flyttar grus en regnig dag.
Flera personer med orange västar går längs järnvägsspåren.
En man i orange väst arbetar med ledningar på en tunnelbana.
En byggnadsarbetare pratar i telefon i en tågtunnel.
Två män i yrkeskläder och hårda hattar samtalar om rapporter.
Två byggnadsarbetare arbetar på en byggnadsställning.
Vit man står på byggnadsställningar med orange jacka målar ett tak.
En arbetare bär en orange väst, hård hatt medan han tickar en byggnad.
Män i orange västar arbetar tillsammans för att lyfta ett föremål.
En man står framför en stor växel.
En byggnadsarbetare i orange väst tittar på en tågtunnel med Kennington-skylt på.
Arbetare arbetar under byggnadsställningar.
En man i orange väst ler när en grupp män jobbar bakom honom.
En arbetare håller en gul maskin på en rulltrappa.
En man i orange overall arbetar under en järnvägsbil.
En man med orange väst bredvid ett tåg arbetar med en handhållen apparat.
Två män bär orange väst med hjälp av en industriell rengöringsmaskin för att rengöra trappor.
Två män med en docka på en rulltrappa.
Män med orange uniformer och falska vingar går nerför en tunnelbanetunnel.
En grupp arbetare på en tågstation.
Arbetare på en ställning håller på att avsluta ett tak i en byggnad.
Två svarta och en vit byggnadsarbetare arbetar utomhus.
Arbetare i orange västar arbetar på tågplattformen.
Byggarbetare lägger tegelstenar i medianen för en tågstation.
En hall är full av stegar och tyg under konstruktionen.
En man som gör underhåll på järnvägsspåren
Män i orange västar arbetar på en byggarbetsplats.
En man som visar hur ett datasystem fungerar.
En flintskallig man med glasögon håller i en gitarr och sjunger in i en mikrofon bredvid sina bandkamrater.
En man spelar instrument och sjunger.
Folk står på parkeringen framför en Central Market.
En flicka kör en leksaksbil medan en ung pojke leker bakom henne
Ett barn i slutet av en slip och glida på en fest
Tre män har ett samtal utanför butiken.
En man i orange kostym svetsar en järnstång.
Orange intjänade män i hårda hattar som arbetar med Jackhammers
Två män verkar ha kul med rullskridskor på trottoaren.
Byggarbete sker på en grusjärnväg.
En Quattro-kran är i drift under tågstationens konstruktion.
En man som står på spåret.
Byggarbetare står på en träbro.
Någon som krigar mot en orange skyddsväst som står på en järnvägsbro.
Fyra män med orange västar och vita hjälmar arbetar på ett järnvägsspår.
Arbetare med orange västar är på en station
Baksidan av en tågarbetare i orange väst och jeans på Kilburn station plattform.
Arbetare i ljusa orange västar på järnvägsplattformen.
En grupp arbetare i orange västar river upp en orange slang i en byggnad.
Nödpersonal med slangar uppradade och nedför trapporna.
En tunnelbanearbetare står bredvid en bil med flera soppåsar inuti.
Byggarbetare reparerar väggar i en tunnelbana.
Byggarbetare som använder sidospår till insidan av en tunnel.
Målare på byggnadsställningar målar insidan av en tunnelbaneterminal.
Många människor i orange jackor arbetar i tunnelbanestationen.
Byggarbetare sliter i ett dike.
Många människor i ljusa orange västar verkar arbeta i en stor byggnad.
En spårvagnsinspektör i orange väst inspekterar spårvagnssätena.
En man som håller i en hatt med orange skjorta tittar på kameran.
En arbetare som läser på ett tunnelbanetåg.
Fyra stadsarbetare med orange västar arbetar på plattformar i en tunnelbana.
Arbetare i orange västar som sätter upp en gul droppduk.
Män i orange västar och vita hårda hattar står på ställningar som arbetar.
Män i uniform som jobbar på en järnväg.
Män står bredvid någon slags hydraulisk maskin.
Byggarbetare står nära spår på natten.
En grupp människor som bär orangea rockar med vita ränder står tillsammans och håller i ett papper.
Under projektets gång samtalade tågarbetare med varandra.
Två medelålders män spelar ett spel i en park en solig dag.
Ett litet barn klappar den lilla vita hunden.
En man jagar en liten flicka i en blommig klänning längs ett asfalterat spår.
Flera människor sitter runt ett picknickbord och dricker öl.
En skara lokala fiskare inspekterar sina nät på stranden.
Föräldrar med små barn sitter vid ett picknickbord.
En ung man håller en liten pojke och ser på honom med kärlek.
En kvinna i röd tröja sitter bredvid en man vid ett bord utanför.
Han ringer sin fru för att säga att han kommer för sent.
En kvinna i en beige jacka som går i en upptagen tunnelbanestation.
Familjen ställer upp för ett foto på ett bröllop.
Tre unga kvinnor och en ung man som sjunger i en hörsal.
En kvinna håller en drink framför ett vitt tält.
En dam tar ett foto med hjälp av en kanonkamera.
Tre kockar lagar mat åt kunderna, en av kockarna är en kvinna.
En grupp barn ser ut som ett stängsel.
En man utan skjorta klättrar upp på en klippvägg med hjälp av ett rött rep.
En flicka i svart tröja häller lite vätska i ett litet glas.
En familj tar en tur på en gul båt.
En grupp människor står utanför på natten och pratar.
En kvinna i röd kostym sitter på ett steg och delar mat med en man i en läderjacka.
En grupp män i gyllene skjortor som sjunger framför en mikrofon.
En man i uniform som bär en låda som går ut från ett flygplans trappsteg.
Tre pojkar på en utomhus basketplan.
En kvinna på stranden sitter under ett paraply.
En man i orange väst har en stor fågel.
Två män står på en sandstrand framför havet.
Byggarbetare arbetar i en tunnel.
Walter Lou Anne Kitty Anställda hejar på framgången med att skapa batteridrivna lokomotiv
En grupp människor som står runt i ett rum.
Här är en bild på en asiatisk kvinna som dricker öl utanför och sitter på en grön bänk.
En kvinna som gör en sandskulptur av en hästs huvud.
En flicka kastar en fotboll på stranden.
Man och kvinna rider cyklar på asfalterad, inhägnad stig nära havet.
Människor går genom en korsning av en stad som består av en grill och pizzeria.
En liten pojke går med en kvinna klädd i rött i rullstol.
Män samlas runt en korg full av färsk fisk när en annan man lyfter den största fisken i luften.
Pops och tjejerna tar 40 blinkningar.
En ung pojke ler längst ner på rutschkanan.
En man knäböjer på marken medan han håller i en banan.
En grupp män i orange skyddsjackor inspekterar motorn på någon sorts spårvagn.
Arbetare i orange overall och strålkastare stående av utrustning.
Två inspektörer i orange västar som kollar ett tågs elektriska dörrar.
Två arbetare städar en byggnad på natten.
En blondhårig man i en blå skjorta omgiven av skärmar som sitter vid ett skrivbord och pratar in i en mikrofon.
En elektriker i en orange overall testar flera kretsar.
En grupp män som bär orangea reflekterande västar och byxor poserar för ett foto.
Pojken är utanför och håller i en sprayburk.
Två unga flickor gör upp och ner muffins former i sanden.
En grupp kvinnor äter på en terrass.
En kvinna i blå skjorta styr sin hund över ett hinder.
En svart och brun hund står på ett tak.
Ett litet barn som bär en röd skjorta som svänger på en fauxdäcksswing.
Ett barn som sminkar en annan kvinna.
En vit hund med krage och koppel är på väg att tugga på en pinne.
Två pojkar skär kött.
En hund plaskar genom vatten och försöker fånga is i munnen.
En man sitter utanför en byggnad.
Silhuetter av män mot en molnig men ändå ljus himmel.
Ett litet barn rider en lila cykel.
En man som bär en vit hatt är mitt uppe i att hamra in en spik i en tjock bräda.
En tjej med röd skjorta springer i gräset.
Barnet i hängslen sitter vid en leksak.
En man och två kvinnor äter mat på en lokal festival.
En svart hund springer på en gård medan en kvinna observerar
En grupp människor som sitter runt ett bord med drinkar.
En grupp människor samlas på stranden, en man bär en surfbräda upp ur vattnet.
Två stora hundar leker i ett rum i ett hus.
En svart hund springer längs stranden.
En grupp cyklister tittar på något på vägen.
En flicka i gul klänning står på trottoaren utanför en affär.
En liten flicka öppnar en födelsedagspresentpåse ivrigt
En dam i blå skjorta och byxor går nerför en lång hall som är glest upplyst.
En kvinna väntar på att få korsa vägen.
En grupp människor i en träningsklass utomhus.
En kvinna klädd i rött är att göra en "rawr" ansikte och en klo imitation med sin hand.
En svart hund går längs gräset och sniffar på marken.
En hund kastar sig över gräset.
Två indianer dansar på ett bröllop med blomblad över hela golvet.
En kille som spelar gitarr på en bänk med en annan man som tittar på honom.
En man som bär jeans, poloskjorta och keps, gaffel i handen, grillar kött utanför på en inhägnad gård.
En man och två barn på stranden.
En brun och vit ko hoppar bort från en svart och vit boskapshund.
En ung flicka klädd för ett bröllop bland brudtärnorna.
En man i smoking och en kvinna i brudklänning lämnar en kyrka.
Två män som spelar gitarr i ett band på en scen.
Närbild av ung pojke med ansiktet och kroppen målade.
Sju byggnadsarbetare som arbetar på en byggnad.
En man i gul jacka som kastar en gul Frisbee.
Man i vit skjorta pratar i telefon medan andra i bakgrunden går förbi.
En grupp indianer sitter i en cirkel och sjunger och slår en trumma.
Ung pojke som cyklar med en äldre man.
Två män sätter upp en stadga och skriver under på ett träd.
En man i en blommig jacka bär hjälm.
En kvinna i svart skjorta svänger väldigt högt på en gunga.
En liten pojke i röd skjorta som pratar på en mobiltelefon.
En man i en marinrock lutar sig in för att kyssa en kvinna i en krämrock.
Det lilla barnet har blå glasögon.
Barnen leker med glittrar på natten.
En blond kvinna i solglasögon som sitter på en bänk.
En brun hund med en liten fotboll i munnen står på en filt
Ett äldre par som tar en promenad tillsammans.
En man i en labbrock som bär glasögon och tittar på en datormonitor.
En ung man i svart skjorta skär kött.
En man verkar förvånad när han blev fotograferad medan han styckade kött i köket.
En man i en cowboyhatt grillar mat på en campingplats barb-que.
Personer av olika raser och etniciteter som väntar på att gå ombord på ett lätt tåg.
En kvinna med en brun jacka sträcker sig in i ett skåp.
2 personer på en strand som begraver en tredje person upp till huvudet i sand.
En kvinna dansar ensam som många människor, i formella kläder, titta på.
Två asiatiska män och en asiatisk kvinna sitter i svarta massagestolar.
En man i ett förkläde grillar majs.
En flicka hängande upp och ner på ett rep över en gräsgräs gräsmatta ovanför en stad.
Den äldre mannen som bär den vita mössan håller upp tummen.
Flera personer lämnar ett kommersiellt jetplan.
En man som sitter på en avsats och äter ett äpple.
Kvinnan i en blå skjorta dricker medan hon lagar mat över en grill.
En man med hästsvans och avskurna shorts hula karvar.
En man i ett rustikt kök lägger mat på disken.
Tre små pojkar står bredvid och på ett staket.
En svart och vit hund går med en blå frisbee i munnen.
En pojke ramlar av sin röda cykel.
Två hundar har båda samma käpp i munnen medan de simmar.
En man som spelar akustisk gitarr framför ett skyltfönster.
En stor brun hund hoppar ner i havet.
Två unga flickor med klänningar och motorhuvar står bredvid ett träd.
En person använder metalltång för att vända en shish kabob vid grillen bland annat grillad mat.
Två hundar står i en pöl och en har en gul tennisboll.
En man som går en hund lägger armen runt axeln på en kvinna med rosa byxor.
Leverans man i en blå baseball keps i en skola.
En pojke klättrar sten i skogen.
Kayaker är i hårt vatten.
Bergsklättraren verkar vara fast mellan en sten och en hård plats.
En motorcykelförare som svänger.
En ung man som spelar elgitarr när han sitter på trottoaren.
En rödhårig kvinna i rosa skjorta försöker gå ner i ett träd.
Ett barn klättrar upp på insidan av ett rött rör i en lekstruktur.
En rödhårig med röd skjorta klättrar upp på trädgrenar.
Vid en liten basebollmatch kallar en umpir "säker" när en spelare korsar hem.
En kvinna i en mönstrad klänning sjunger in i en mikrofon.
En grupp människor på mobiler som tittar på himlen.
En flicka håller i ett rep ovanför vattnet.
En man i ett laboratorium häller en klar vätska i en maskin.
En man i rutig kostym som skakar någons hand.
En svart och brun hund springer på stranden.
Tre barn spelar fotboll i sanden.
En flicka tittar över en pojkes axel när han läser en bok.
En kvinna i blå byxor är bergsklättring.
En liten pojke i badrock sitter i en metallstol.
En kvinna i blå sweatpants lutar sig mot sin ryggsäck i skogen.
En kvinna med vitt hår mejslar på en ofullbordad skulptur.
En ung pojke lutade sig framåt i ett barns sving.
En grupp människor som spelar ett spel med en tennisboll på en strand.
Två hundar springer genom gräset bredvid en gata.
En brun hund som springer i fält av långt grönt gräs.
En liten ligapojke som gör en träff.
En ung, vänsterhänt smet i baseball ögonblick efter att han gjorde en träff med en catcher i närheten och en publik i bakgrunden.
Lilla flicka som håller på att svalna i poolen.
En ung flicka med glasögon sitter och håller två amerikanska flaggor.
Barn i hjälmar spelar hockey utomhus.
Två män i baseball hattar säljer sparris och andra grönsaker från en utomhus monter till en kvinna som bär en grön väska.
En brun hund hoppar genom ett fält.
En man i en nummer 11 skjorta redo att spela fotboll på fotbollsplanen med tusentals människor tittar på.
Det finns många människor som bär hjälmar som rider på cyklar.
En man i orange skyddsväst går mot vissa byggnader.
Tre hundar tävlar vilt runt en kapplöpningsbana.
Ung man klädd i svart med vita tennisskor, liggande på en stor grå sten.
Mörkfärgad Mercury bil parkerad framför PNC Bank.
En ung flicka i simglasögon gör ryggsim i en pool.
En ung pojke i gul skjorta som går på stranden och bär en surfbräda
Tre drakar är i luften framför en bergskedja.
En flicka övar sin tjänst på parkeringen.
Fyra kvinnor i liknande röda kläder sjunger och använder trummor som de utför.
Farmer säljer konserver från en skåpbil.
Närbild av hund i profil med munnen öppen.
Två barn låg i gräset.
Folk tittar på kläder och andra föremål på en utomhusmarknad.
En svart hund som står i vattnet.
En person med badmössa och glasögon tar ett andetag.
Fem män står i en båt.
En ung barfota flicka hoppar upp i luften medan hon spelar leksaksgitarr.
En man som leker med en bollleksak med sin bruna hund.
En kvinna klädd i svartvitt röker en cigarett i ett gräsbevuxen område.
En svart hund dränkt i flytande hoppande till gräset.
En flicka studsar i en sele med en byggnad i bakgrunden.
Barnet sitter på sandstranden.
En man med huvtröja och jacka sitter på en bänk i en park.
Två hundar går längs grusvägen.
En pojke i en orange "Spring Hill" boll lag uniform, pitching bollen.
En pojke i en pool som bär Spiderman-floaties.
En kvinna som leker med lekredskap medan ett barn tittar på.
En asiatisk man som sitter på en stadsgata.
Flera människor står och sitter på ett gräsfält och ser en hund hoppa över en man för att fånga en apelsinfrisbee.
En brun och vit hund springer över gräset.
En man i denimshorts och en halmhatt fiskar bort från klipporna.
En kampsport klass äger rum i Ourense, Spanien.
En ung pojke och flicka sover i en säng.
En liten pojke sitter på betongväggen vid havet.
En man i en rishatt bär många föremål.
Simlärare visar unga flickor hur man flyter.
Fyra kvinnor i röda baddräkter uppträder i vattnet när en skara människor tittar på.
En liten pojke i Hawaiis shorts spelar i en sprinkler.
En kille i svart läder motorcykel kostym en hjälm på en silver motorcykel.
En skara människor njuter av solskenet på en plaza.
En kvinna pressar en man i rullstol; i bakgrunden är en båge.
Folk går genom en fullsatt gata.
En ung pojke leker i fontänerna och skjuter upp från marken.
Två hundar springer i vattnet.
Ett barn håller i en kopp och leker med en leksaksvattningsburk.
En liten hund leker i gräset.
En vithårig man lägger ner sin käpp och hatt och vilar bredvid ett träd.
Den upphängda målaren målar en vägg.
En grupp unga tonåringar försöker fånga ett föremål i en utomhusgränd.
Tre män utanför på uteplatsen i en byggnad.
En flicka knäböjer på en rund fontän som sprutar vatten i luften.
En ung pojke klättrar upp på klippväggen.
De tre svarta hundarna simmar mycket nära varandra.
En man tittar över ett räcke i vattnet.
En ung flicka som jagar bubblor medan hon springer på en trottoar av skiffersten.
Ett lyckligt ungt par som har ett glas gnäll och pratar.
Två damer som sitter vid ett bord har ett skratt.
Kvinnor håller upp två karikatyr porträtt av sig själv under middagen.
En person klädd i allt blått går nerför en väg med höga träd på vardera sidan.
En man som ritar en bild av två kvinnor.
En man med en handskada går med en käpp i en park.
Två hundar möter varandra i ett fält
En man i grön skjorta står mellan två bilar som håller upp 3 fingrar.
Kaukasisk kvinna i svart klänning, nära ett gammalt trästaket.
Två kvinnliga tävlande går ut med sina hundar i en hundshow.
En cementbil häller cement på gatan.
Ett barn, som sitter vid ett bord, håller en smörgås i sina händer och gråter.
Folk som sitter eller står på en buss.
En medelålders gift kille i gul skjorta svettas och spelar en brun gitarr
En löpare jagas av en man i en pingvindräkt.
Två hundar springer genom grunt vatten i en vik.
En stor, röd traktor drar en platta längs en grusväg.
Det finns en stor grupp människor som står i gräset och de flesta av dem håller händerna i luften.
En man som springer barfota på gräset.
De två grå hundarna försöker få ett rött föremål.
En förbipasserande och en byggarbetare på trottoaren.
En kvinna som bär shorts håller ett barn bland en skara av mestadels barn utanför i en stor fontän.
Två asiatiska tjejer uppträder i kostymer.
En kvinna cyklar genom en upptagen marknadsplats.
En man lyfts av en annan man i en asiatisk kampsport rörelse.
Två pojkar med baseballmössor sticker ut gröna färgade tungor.
Två hundar skäller bakom ett stängsel.
Ett litet barn springer nerför en grusväg täckt med döda löv.
En man är i en frisörs butik och klipper sig.
En man står bredvid en stor, färgglad fågelbur som innehåller fåglar.
Två afroamerikanska barn läste en bok.
Tre personer står i en gång mellan två hyllor staplade med böcker.
En blond kvinna som försöker ha klackar i en skoaffär.
En vit kvinna sitter och läser medan hon är omgiven av sex små svarta barn.
Byggnad med svarta som sitter utanför i ett land i tredje världen.
En kvinna i grön skjorta som står på ett podi.
En kvinna med brunt hår ler och bär ett konventmärke.
En kvinna i svart kostym står och ler framför en annan kvinna i röd jacka.
En grupp vandrare tittar på en butiksdisplay.
En man med en gul skjorta som står bakom ett svart podi.
Laura Bush talar vid en konferens om global läs- och skrivkunnighet.
Kvinnor i afrikansk dräkt sitter utanför medan en i väst går förbi.
Afrikanska amerikaner sitter på stolar i ett klassrum.
En man pratar medan två människor är nära honom.
Tolv barn sitter på marken.
Det är många barn som har kul på en fest.
En ung flicka städar marken med en trasa.
En mamma sitter ute på en stol medan hon håller sin dotter i knät.
Ett barn i en sving.
En ung afroamerikansk pojke som sitter på en träbänk i ett bibliotek och tittar igenom en bok.
De skriver medan de bär blått.
Tre hundar springer bort från en fläck av icke gräsbevuxen yta och lämnar varandra bakom sig.
En man och en kvinna som möter varandra på en bänk.
Två bruna soffor vänd mot varandra över ett soffbord fullt med tidningar och tidskrifter.
Människor går på grusväg med två lastbilar
En man i blå skjorta och en kvinna i rosa kjol sitter runt andra människor i bakgrunden.
En grupp människor sitter i skuggan under ett träd.
Två män i uniform håller upp skylt med små barn.
En ung flicka i blått hoppar upp i luften.
En vit hund springer nerför en stig mellan buskarna.
Hunden går i det grunda vattnet.
En gråhårig man med glasögon sitter på en stor bänk med benen utsträckta.
En stor kvinna står på gatan.
Kvinnan i rosa går en promenad genom ett fält.
En man i en quiltad jacka sedd bakifrån står framför en korgstol.
Sex unga pojkar, en afroamerikan, en latino och de andra kaukasiska, står framför ett staket som bär olika typer av kläder, och fem av dem håller sina öron.
Två tvillinghanar viker ihop en blå handduk.
En grupp män som sitter på golvet i ett fönsterlöst rum.
Små pojkar i sporttröjor leker med en gul boll.
En ung man rakar av sig skägget med rakskum och rakhyvel.
Flera människor sitter inne i ett mörkt konstgalleri.
En professionell idrottsman kliver fram till plattan för att göra en sväng på bollen.
Två hundar leker med en käpp i vattnet.
En man i gul skjorta och khaki shorts balanserar på en metallkedja.
En man fyller upp en gammal hink med sand.
Ett litet barn i en ljusblå overall sitter högst upp på ett rött plastglas.
Steers och man njuter av en dag på stranden.
Infödingen fiskar i en utgrävd kanot på en blå grön vik.
En man spelar munspel i en restaurang som står framför dig.
En man med många tatueringar och kroppsgenomborrningar sväljer ett svärd i en föreställning på en utomhusfestival.
En man blandar något i en mycket stor skål.
En man i randig skjorta spelar gitarr för flera människor som står runt honom.
En kvinna som bär en hink med blommor.
En man, som bär en blå skjorta, bär hörlurar och arbetar med ljudutrustning.
En polis tittar på en annons i ett fönster
En pojke i blå fotbollströja och shorts står och ser två andra barn spela fotboll.
En liten flicka i rosa skjorta som ska gråta
En mountain bikeer i rött rider på en skogsstig.
Fyra personer tittar genom ett stängsel.
Cowboy i blå och röda byxor blir bortkastad från en häst.
En vit hund som springer genom gräset.
En kvinna är utanför och tittar över havet när solen går ner.
Mannen tävlar sin cykel nerför kullen.
Ett lyckligt gaypar som tar en promenad genom en park.
Fem asiater sitter runt ett runt bord.
Folk hänger upp och ner när en berg-och dalbana utför en spiralslinga.
En kvinna håller en linje på en segelbåt.
Hunden hoppar genom vattnet.
Möbler inuti och utanför en flyttbar lastbil.
Ett litet barn i en Izod-skjorta håller en mobiltelefon i örat.
Soldaten sitter ovanpå jeepen och håller ett kulsprutor och en soldat som sitter inne.
En grupp på fem poliser på motorcyklar rider på en stadsgata.
En pojke som bär födelsedagshatt spelar i en pöl.
En fotbollsspelare som springer med bollen under en match.
En man reparerar en segelflygplan på en solig dag.
Fyra män utför arbete i en smuts mycket, nära en byggnad, med hjälp av en soptipp.
En person i orange hjälm åker skateboard på en ramp.
En man i brun skjorta håller en blå hatt över huvudet och en röd hatt på armbågen.
En utomhusfestival verkar äga rum.
En yngre man med glasögon sitter på en gräsplätt bredvid andra människor.
Den här ungen säger att bergsklättringen är en kick!
En man i en tvivelaktig botten hjul sin livsmedelsvagn över en samling på gatan.
En man som sitter på huk i en park och tittar på något i fjärran.
En grupp människor som är nakna och rider cyklar på gatorna.
En vit man på en telefon sitter vid ett mycket rörigt skrivbord.
En man i en röd knapp-down skjorta undervisar en klass i ett klassrum med blå målade väggar.
En lärare fixar en liten elevs hår.
En pojke med blå hjälm och grå byxor kliar.
Två byggnadsarbetare bär hattar och orange västar.
Byggarbetare klädda i skyddsvästar och hattar inspekterar sitt arbete.
En man som står bredvid ett fortkörningståg och tittar på sin mobil.
En ung man sparkar en fotbollsboll i ett tomt tegelområde.
En man som spelar boll vid solnedgången.
En liten hund skäller på en brun och vit ko.
En grupp män står utanför ett pizzaställe.
En liten hund hoppar upp för att möta en gul fotboll.
En man i blå och gula shorts håller handen över vatten.
En kvinna som bär en vit bikini övredel får hjälp av en man att korsa en vidd av vatten.
Tre personer sitter i ett rum med cykel och skoter.
En kvinna i förkläde håller en fisk och det finns en blå gryta och flera andra ingredienser på bordet.
Ett barn står framför en dansande bröllopsfest.
Medan en man i röd tröja sitter på en bänk samtalar han med en man i en lila kofta.
En brun hund hoppar högt i gräset.
Det finns en person som står på en trappa utanför en Costco-butik.
En grupp bilar parkerade på en kulle
Två män på en konsert skriker.
En hund vadar genom djupt vatten medan han håller i en pinne.
Två män med orangea skjortor som knuffar barn i barnvagnar under maraton.
En liten pojke blåser bubblor genom ett trollspö som hans mor håller i.
En ung flicka och två unga pojkar som leker med scooters på en docka under dagen.
En ung flicka i rosa och vit klänning kramar en examen.
På det här fotot står en ung pojke klädd som en basebollfångare på knä bakom hemmaplan.
En liten pojke rider en gul cykel över ett torg.
En svart hund håller en svart fågel i munnen.
En kvinna i grön klänning väntar med sitt bagage.
En man som ligger på ett sittansikte och kanske sover.
En ridsport hoppar upp i luften på hästgården.
En brun hund blir blöt i vattnet.
Tre unga pojkar blinkar med händerna och ler.
Två män och en dam går längs en landsväg med öl, apelsinjuice och elektronisk utrustning.
En del människor äter på en matplats.
En liten flicka i vit klänning och inga skor går längs en grusväg i Amerika.
En vuxen drar ut ett barn ur en bollhåla.
Mannen kastar en tennisboll för den bruna hunden att hämta.
Folk rider cyklonen spänning rida på Coney Island nöjespark.
En ung flicka i rosa skjorta håller i ett par hörlurar.
Tjejen väntar på att bollen ska komma ner när hon spelar tennis.
Två pojkar leker med en hulahoop på gården.
En ung man sitter på vägkanten med sina tillhörigheter.
En man och en kvinna sitter med en skylt och läser "Det är en fin dag för ett gaybröllop."
En liten pojke tar en bild i parken.
En svart man i vit kostym och hatt håller i en pappersmugg.
Två hundar springer mot varandra över sanden.
Två flickor är i ett säcklopp.
Tre kvinnor står nära en upptagen korsning.
En svart och vit hund ser tillbaka när han går på stranden.
En europeisk bonde lägger ner hö för att hindra floden från att erodera.
Två grupper av människor sitter i ett bås i en middag.
Tre kvinnor hoppar samtidigt av en kuststad.
En liten flicka som håller en frilly vit klänning ut för den andra lilla flickan att undersöka.
Folk tittar på TV medan de äter.
En ung flicka framför ett bibliotek springer genom en fontän.
Den vackra unga flickan går genom röret.
En hunds huvud ligger i knät på en person som äter av en liten tallrik.
En pojke och flicka leker i en pool.
En brun och svart hund som går på stranden
En man i vit keps och skjorta handpallar en liten blå båt.
Ett leende barn håller ett långt gult och grönt objekt medan man tittar på ett annat barn som håller ett liknande objekt.
En liten pojke i baseballkläder som svingar ett slagträ.
Ett barn med glasögon och en badmössa som simmar i en pool.
Unga pojkar tränar simning i en inomhuspool.
Barn i blå klänning som håller sandal i ena handen och äter blått bomullsgodis med andra handen.
Ett band som spelar på scen för en massa människor.
En flicka i rosa skjorta och en man i vit skjorta går på ett fält.
En mindre vit hund och en stor herde som leker nära två personer.
En man med dreadlocks, promenerar längs en gata café medan strimla en gitarr
En tonårspojke utför ett trick med sin skateboard.
En man i grå skjorta står framför ett stativ med skålar med färgglada puder.
En kvinna i lila ridande uniform rider en häst genom ett fält.
Unga pojkar med ryggsäckar går nerför gatan förbi en stor byst Buddha
Familjen kopplar av i gräsmattan stolar och dricker.
En liten pojke med ett smutsigt ansikte ligger på en färgglad matta.
En konstnär som väntar på att teckna en person på gatan.
En grupp unga pojkar som stod nära en annan pojke som satt på en gunga på en lekplats.
Två kvinnor i vita klänningar promenerar genom en park.
En man med en cigarett och en kvinna i en blå skjorta kysser i en bar.
Två män med orange väst lutande över ett räcke.
En hund hoppar på ett fält medan en annan hund står bredvid det.
En kvinna i röd skjorta står framför en komålning.
Ett svart labb hoppar från en brygga ner i en damm.
En monter med många olika torra livsmedel, såsom nötter.
En familj äter vid ett bord och dricker vin, med två barn, modern, fadern och en oidentifierad kvinna.
Folk pratar vid ett evenemang i en park.
En grupp människor samlas runt picknickbord i en park kantad av träd.
Ute i en park står åtta personer nära ett skräpigt picknickbord.
En grupp människor på en livlig gata.
Kvinna i rutig skjorta och kjol håller växt och leende.
En flicka med rosa hatt går bredvid ett får på en dammig stig.
Två pojkar står och surfar.
Ett litet barn tycker om att spela i en bil som har den tecknade karaktären "Barney".
En liten flicka med blont hår som tittar på publiken.
En man som knäböjer vid en ljusröd kajak med flera kajak- och kanotskyltar bakom sig.
En brun hund och ett svart hundslagsmål.
En gammal kvinna i en möbelaffär, en liten hund tittar på när hon går sin väg.
En man på en surfbräda som rider på en jättevåg.
Den unge pojken fladdrar lera vid barfotaflickan i dammen.
En man håller en turkisk flagga utanför fönstret på en bil.
En man i blå skjorta och brun baseballhatt äter ägg på en restaurang.
Pojken glider nerför rutschkanan med utsträckta armar.
En man i neongrönt städar upp utanför en byggnad med lite graffiti.
En liten pojke poserar på en stenvägg utanför.
En liten grisstjärtad flicka i en rosa tröja tar tag i en ung pojkes ben.
En ung pojke och flicka som leker.
En hund biter en katt medan de ligger på en säng tillsammans.
Det finns sex arbetare på en byggarbetsplats.
En pojke sitter vid ett bord och skriver i sin anteckningsbok.
En far och hans barn sitter på en bänk vid en grill.
En tennisspelare bär en röd skjorta på väg att slå en tennisboll med sin racket.
En kvinna som bär vit skjorta håller upp en limpa bröd.
Två tjejer med långt hår som hoppar på en studsmatta.
En kvinna med blommande lei spelar gitarr.
En man med mustasch och svart hatt håller ett litet gult föremål upp till kameran.
Två svarta hundar simmar i en pool.
En flicka som använder en rosa penna för att anteckna ur sin bok.
Ung vuxen i grön skjorta med rödhårig skrift på ett papper.
En ung pojke blåser bubblor på en gräsbevuxen gräsmatta.
En man med grönt pannband arbetar på ett byggprojekt.
En kvinna i grön bikini ligger i vattnet.
Folk är upptagna med att äta på hotellet.
Flera människor är i ett rum stirrar på en vägg med projicerade bilder på den
Flera personer spelar instrument i ett rum tillsammans.
En pojke knuffar en kundvagn med en annan mindre pojke stående upp i den.
Ett barn snurrar en handhelikopter i ett gräsfält.
En ung flicka tittar på alla färska produkter som finns på marknaden.
En röd hund står i en stenig strand, dess fötter i havet.
Två hundar står bröst djupt i vatten, bredvid en pinne.
En stor brun hund och en stor svart och vit hund som springer tillsammans
Två bruna hundar leker i grunt vatten
En informellt klädd orkester repeterar i en tom hörsal.
En ung kvinna i en tanktopp och culottes bär på ett barn.
Barnet håller en kamera på nära håll.
En man knuffar en barnvagn nerför en våt väg med ett barn som går längs sidan.
En man sitter ner medan han svetsar ett föremål.
En familj hoppar in i en sprängflotte i sitt vardagsrum.
Det svarta och vita djuret är i gräset.
En man i röd skjorta på gatan gör ett brandtrick.
En grupp musiker samlas för att spela musik.
Två nakna kvinnor målade svart och vitt rider cyklar på vägen.
En topless kvinna är täckt av lera.
En man en blå skjorta matlagning mat på en grill.
En afrikansk kvinna som stod nära ett staket vid vägkanten.
En man med rutig skjorta och grön hatt klipper gräsmattan nära trottoaren.
Ett par i en restaurang håller hand.
En orientalisk kvinna som bär hatt går nerför den livliga gatan.
En hund med frisbee som badar i en sjö.
En svart hund och brun hund springer runt i sanden.
En grupp barn hoppar in i en pool.
En kvinna i brun kostym och luddiga svarta vingar cyklar
En man spelar tangentbord med en annan man som spelar trummor.
Pojkar står utanför ett tegelhus och en pojke börjar springa.
En upptagen kvinna poserar snabbt för en bild medan moppa köket.
En grupp barn står under några banderoller och sträcker armarna över huvudet.
En äldre man som går nerför gatan otrygg på människorna omkring honom.
En pojke i vit t-shirt plaskar i grunt vatten.
En bil står parkerad på en graffitifylld gata.
En ung, blond flicka i en fe utstyrsel rider en rosa och lila trehjuling.
En grupp barn springer med en hund nerför en gräsbevuxen kulle.
En liten pojke med blondin leker med sand och en spade.
Två män utan skjortor tvättar ett tak.
Två personer går längs stranden vid solnedgången och varnar en grupp människor.
En tennisspelare i en vit outfit träffar en tennisboll.
En man som ser ledsen ut när han håller en näsduk på en stadsbuss.
Två killar är inhägnade i ett jordområde.
En ensam swinger på en svängtur på marknaden.
Två män som bär på fiskestänger som går längs stranden.
En man i vit skjorta med glas som rör om i maten på spisen.
Två kvinnor tar utomhusfotografier på en askbana.
Två bruna och vita hundar, en hoppar över en stock medan den bakom springer genom gräset.
En man tar av sig skorna, sitter på bänken och tittar på den stora fontänen.
En man och en kvinna i svart sitter vid köksdisken och tittar på en kvinna i en röd tanktopp blandar deg på en skärbräda.
Folk går nerför en trottoar på en strand.
Tre kvinnor är i olika poser på en stig kantad av bambuträd.
En man i svart skjorta läser på sidan av en skål.
En dam i ett kök står framför spisen och steker något i en stekpanna.
En pojke som går genom stolar och bord på Au Bon Pain.
En man i denim overall rider en Segway nerför en strandpromenad.
En vuxen som håller i ett mycket litet barns ben medan han sitter i en hängmatta.
Tre kvinnor solar på en stenformation som gränsar till en vattenförekomst.
Mannen utför stunt, damen bryter block på magen med slam hammare.
Två vita hundar springer sida vid sida i grönt gräs.
Två män jobbar på en stålstruktur.
En stor grupp människor deltar i ett maraton längs en stadsgata.
En grupp hejaklacksledare i svart och orange kläder hejar på.
En man i blå jacka är uppe på en stege som får hjälp av en kvinna i en röd jacka
Två män i en bygghatt och reflekterande skyddsvästar på jobbet.
En gymnast böjer sig över på en gul matta på gräset.
Barn spelar i en fotbollsmatch.
Flera kvinnor, klädda i rosa "Energizer" kaninöron, pekar åt höger.
En svart hund som hoppar från en docka i vatten.
Fiskare arbetar sina nät närmare stranden medan en båt sitter i vattnet som är anslutet till näten.
Stor hund och katt stirrar på varandra på en tegelsten.
En man går på stranden och lämnar några fotspår bakom sig
Ett barn sitter på ett däck och håller en leksak.
Klippor omger en äventyrares fötter och gräver sig ner i en underjordisk grotta.
En gammal man sitter på en bänk med utsikt över vattnet.
En glassbilsanställd sitter på sidan av glassbilen.
En publik hänger framför en rosa "finish" sinus.
Ett ungt barn leker med sina plastleksaker på trottoaren, medan en kvinna med en shoppingväska lutar sig mot en grön metall bar.
En kvinna och två barn med hatt går nerför ett spår.
En vacker dam sitter vid ett bord klädd i en ljusblå klänning.
Folk samlas för något evenemang i staden.
Den lilla vita och bruna hunden simmar i en pool.
Unga flicka poserar med publik i bakgrunden
En pojke i röd väst och vit karatedräkt sparrar med en pojke i blå väst.
Tre brudtärnor i blå klänningar håller tåget till brudens bröllopsklänning.
En kvinna i brudklänning inspekterar en bukett.
Brudtärnor och brudgummar poserar för ett foto med paret att gifta sig.
Ett gift par poserar för bilder på en gräsbevuxen bergssluttning en molnig dag.
Ett gift par som ser ut vid vattnet.
Två personer sitter i mörkret nära en flammande eld.
En kvinna springer i ett maraton.
En eventuellt berusad man ligger på marken bredvid en livlig väg.
En äldre man har ett litet spädbarn som är inlindat i en blå och vit filt.
En man i parken som klättrar lite.
En ung kvinna, topless förutom färg eller lera.
En skateboardåkare gör ett trick i luften på en skridskor ramp.
Två hundar som leker på en skolgård
Vid ett tegelgolv nära stranden sitter en medelålders vit man omgiven av en vit familj och målar ett porträtt av någon.
En grupp barn får lära sig att använda datorer.
Vi svär trohet till vad du vill om du bara ger oss lite mat.
En kvinna med en rosa skjorta som målar en stjärna på den amerikanska flaggan.
En hemlös man i vit mössa står bakom stora, orangekottar.
Två flickor som sitter på marken
Människor som bor i slumområden visar hur de försöker städa.
Två pojkar som står i ett fattigt område ovanpå en sophög.
Den ene sover, den andre hoppar på sin säng, båda bär vitt och ser ut att vara på indisk härkomst.
En liten pojke och fyra kalkoner som går
Flickan svänger glatt på en sväng utanför.
Skateboarder utför ett spektakulärt trapphopp.
En byggnadsarbetare bär två och fyra, framför en nybyggd trävägg.
En man går med en ko nerför en grusväg.
En hawaiiansk man utan skjorta på sig och bär en rosa blomma i håret och en grön wrap spelar ett instrument.
En färgstark parad till ära av bilder avbildade på en tavla.
I ett vardagsrum förbereder sig en ung pojke som bär ett leksaksstetoskop för att lyssna på en kvinnas hjärtslag.
En flicka som sträcker sig ner i vattnet medan hon står vid kanten av en flod.
En kvinna med lockigt hår tittar genom en stor uppvisning av plånböcker på ett bord.
En hund jagar en hjort in i skogen.
En man som bär en blå rutig skjorta biter i lite mat.
En asiatisk man som borstar tänderna vid ett vitt handfat.
En flicka svingar en ung pojke nära en välvd dörröppning.
Ett lyckligt barn bär en orange livväst.
Två hundar springer i ett fält av högt gräs.
En grupp människor som sitter på en soffa och dricker drinkar.
En mor och dotter går på gatan och passerar en man som läser en tidning.
Nummer fyra hunden framför andra hundar.
En man i svart jacka med vit rand nerför ärmen ler.
Två damer sitter och tittar på något.
En välklädd man sover framför ett skyltfönster och annonserar böcker.
Sittande ungdomar försöker följa instruktioner och slutföra en modell
En person på en motorcykel som slår en wheelie i en parkering.
En liten hund jagar en tennisboll på trottoaren.
En kvinna visar en hund med mycket långt hår på en hundshow.
En man med vitt hår, blå jeans och en vit T-shirt som skär ett objekt.
Två män interagerar med någon sorts mekanisk apparat som är monterad på en vägg.
En indisk man med en stor mobiltelefon.
En barfota kvinna med en tanktopp som tittar på leksaker i en gång i en affär.
En färgglad klänning person poserar med ett blått och vitt paraply.
En man svetsar utan ordentlig säkerhetsutrustning på.
En liten flicka tar en bild utanför.
Kayaker i skyddande hjälm och blå kajak håller sig flytande i rasande vatten.
En person som hoppar från en hög klippa.
En man i ateljén tittar på sin pågående skulptur.
En pojke svänger i luften.
En brun och vit hund går bredvid en man på en skateboard.
En arbetare tittar ut i fjärran medan en China Shipping låda sitter bakom honom.
Den grå hunden blundar.
En ung pojke rider en röd häst.
En liten hund tittar på en tennisboll i luften och en papegoja sitter i närheten.
Ett blond barn går förbi ett skyltfönster.
Två äldre män utanför lastning eller lossning av en släpvagn full av stora vita cylindrar.
En vit hund sitter på en stenig gräsmatta.
En liten pojke i shorts och en röd skjorta, luftburen på en uppblåsbar rutschkana.
Polisen på motorcyklar eskorterar en bilkortege.
Två män pratar, yngre och äldre, medan den visa gamla ugglan lyssnar, i tystnad.
En man med solglasögon sätter ett chip i munnen.
Två män hälsar varandra med en kram.
Folk rider skotrar genom en fullsatt gata.
En flicka i rosa hatt tittar ut över en vattenpöl.
Den lille pojken böjer sig ner för att titta på ett djur.
Flera ungdomar i svarta och vita skjortor och blå jeans går nerför en gata.
En svart hund jagar en röd boll genom vattnet.
En kvinna stryker kläder i ett sovrum med trägolv.
En man i en folkskara höjer sina armar på bön.
En grupp människor samlades runt en tegelbyggnad som har tre män på sig.
En ung flicka i lila baddräkt som tar en paus vid poolen.
En svart man köper nåt i kassan i en affär.
En ung man tänder en tändare medan en annan tittar på.
Två män kramas i en folkmassa framför en tegelvägg.
En softball spelare springer mot hemmaplattan.
En liten grupp arbetare verkar arbeta på gatuutgrävningar eller reparationer medan en kvinna och en man går förbi dem när en svart sedan kör förbi.
Byggarbetare häller betong för att fylla ett hål på sidan av vägen.
Två män arbetar med en cementblandare och häller cement i ett hål på en gata.
Personen på cykeln bär rött.
En äldre pojke med armen runt en yngre unge under ett sequoiaträd.
En man som gör ballongfigurer under ett utomhusevenemang.
Ett litet barn och ett barn leker i slutet av en rutschkana.
En man med buskigt skägg och rosa skjorta ler.
En kvinna tittar på taket medan hon tar av sig hatten.
Ras hundar mitt i luften medan de springer.
Två pojkar klädda i vita kåpor som springer på en stig i ett fält.
En gammal man står framför en rasande byggnad.
En man med ryggsäck sitter på en fallen stock vid floden.
Två personer står med en naken gitarrist på en livlig gata.
Tre killar jobbar med en stor glasram.
En hund med en pinne följer en annan hund genom vattnet.
Är äldre kvinna i en svart topp uppmärksamt läsa en bok vid köksbordet.
En leende pojke flyter i en pool.
En stor brun hund simmar mot kameran.
En man och kvinnor sitter på en strand medan solen går ner.
Den unga damen med den röda skjortan är framför publiken.
Tre polisbilar behövs för att gripa en misstänkt.
En skolgrabb som sitter på en citronjuiceaffär känner att han vill smaka på den där saften.
En leende kvinna håller en tårta nära en man.
Medan andra ser på hoppar en ung flicka ner i en bassäng när en kvinna sträcker sig efter henne.
Urban Tree arbetare beskärning ett träd medan upphängda av en sele.
Män som sjunger blues i en av de vackra orkesteravsnitten tack vare Shell Corporation of America.
Ett barn med huvudet avskuren från en ko.
En hund hämtar en tennisboll i en patch av grönt gräs.
En hund sträcker sig över det gröna gräset.
En asiatisk flickas vatten växer bredvid uppfarten när en dam går förbi på trottoaren.
Den lilla ungen svänger i trädgården.
En brun och svart attackhund tränas av en man som håller i en pinne
Den stora beige hunden springer genom gräset.
En kvinna, i den rosa skjortan, spelar Jenga, medan två unga vuxna tittar på.
En hund hoppar över ett hinderbana stängsel.
En flicka i en blommig klänning gråter på en sanddyn.
En man har utsikt över ett stort, snöigt berg.
Två personer som bär jackor går förbi en museiutställning medan flera människor omger utställningen.
En ung flicka i rosa byxor vatten krukväxter.
En skara människor har samlats bredvid ett fält av färgglada vilda blommor.
En snabblöpande Greyhound under ett lopp.
En orange kanot riktad mot två andra kanoter på en sjö.
En kvinna som tränar kampsport i ett gym.
Damen som bär halmhatt och flip-flops ser det kastade föremålet flyga genom luften.
Tre kvinnor och en liten flicka leker med en liten valp.
En liten pojke i grön skjorta håller i en stor orm.
En flicka som sitter på en vägg nära vita kors i marken.
En man i gul jacka rider en gul cykel lastad med flera paket på gatan.
Fem små flickor i gult spel i ett rum med leksaker.
En kvinna som bär en svart sjal går ut ur en byggnad.
Ett barn med en tröja håller en penna i munnen.
En pojke i blått dricka från en kopp med andra barn i bakgrunden.
En kogård vid foten av ett berg nära en sjö.
Tre kajakpaddlare färdas i vattnet längs snötäckta berg.
Barn spelar ett tv-spel tillsammans.
En pojkfångare i hjälm som sträcker ut sin handske för en fångst.
En man står och tittar i fjärran när solen når toppen bakom en trästruktur.
Ett par sitter på en klippa med utsikt över en dal fylld med träd
En kvinna i en huvudduk i öknen
En liten flicka i rosa baddräkt skrattar vid en pool.
En brun hund bredvid en stenbänk.
En grupp människor klädda i karateuniformer sparkar alla upp i luften.
Två hundar leker bogserbåt med en skiva, i knähögt vatten.
En man och en kvinna står under en tegelbåge och läser tidningar.
En man i England och en jersey står på ett gräsfält.
Ett barn som står hukat på en trädlem.
En man går in i skuggorna av en passage.
En hund simmar genom vattnet och håller en käpp i munnen.
En byggnadsarbetare står högst upp i en träkonstruktion.
De här männen är instängda och bygger vad som ser ut som en stiftelse.
Ett barn hoppar upp och ner på en studsmatta.
Ett barn i vit klänning passerar ett bord bredvid en damm.
En person rider på ett djur framför en folkmassa.
Två kvinnliga artister som bär kostymer står på gatan bredvid en byggnad.
Ett barn som bär hatt och en vit skjorta sitter.
Unge pojke som lagar mat i en grill på bakgården.
En man hoppar i luften på en snötäckt bergssluttning.
Fyra honor, varav ett barn med mask i rosa skjorta.
En ung pojke verkar ha roligt i en park.
Två män står vid mitten av en stadsväg.
En publik tittar på löpare under ett maraton.
Två killar står utanför en byggnad som har sprejmålats med ord.
En liten pojke skateboards på en cement ramp.
En brun hund som skakar av sig vattnet
En gråhårig man står i vattnet med en gul hink.
En kvinna som bär en halsduk på huvudet sitter bredvid en ung pojke i blått.
Två hundar tittar upp på en person.
En liten pojke i röd skjorta och baseballhatt knäböjer i grunt vatten med en gul hink full av sand.
Två små hundar jagar en röd randig boll.
Ett barn sitter ovanpå en stor stubbe.
En liten pojke som äter en röd isglass.
Medlemmar i ett band uppträder klädda i vitt medan trummisen sitter bakom dem.
En man står på gatan under kvällen.
En hane och två honvandrare ställer sig framför ett bergigt landskap.
Det finns ett litet barn som leker på en lekplats.
En grupp människor sitter nära havet.
Två små barn, en pojke och en flicka, stod nära en gatuförsäljare och pratade.
En brun hund som känner lukten av en grå hunds svans.
En kvinna i bröllopsklänning borstar tänderna.
En fotograf kikar ut mellan klippiga kullar för att ta en bild.
Person i rosa skidor bär skidor på en sluttning.
Solen går ner bakom en bro medan en man cyklar.
Flera människor går längs en naturskön enkelriktad motorväg.
Ett litet barn sitter på några kuddar med en grön bricka med hackad mat framför sig.
En svart och vit hund går genom ett fält.
En flicka med kortklippt hår lagar mat på en grill.
En pojke ser sur ut när hans far tittar på kameran.
Svart hund med svart och brunt ansikte som rinner genom vatten.
En militärmedlem talar med en annan medan han är ute på gatorna.
En man med skrynkligt skägg passerar ut flygblad nära några cyklar fastkedjade vid en grind.
Flickan håller i en grön boll.
En asiatisk flicka som bär på en rosa väska går sin väg nerför en livlig stadsgata.
Unge man visar upp sig genom att dyka från en klippa framför sin tjej.
De två små hundarna springer genom gräset.
En kvinna med vit skjorta som går nerför trottoaren.
Kvinnan bär svart solhatt, svart klänning och svarta Ugg-täppor, som går på ett torg.
Två unga pojkar i kostym brottas.
En asiatisk man och kvinna möter varandra och gör arga ansikten.
Två kvinnor går över en gata tillsammans.
Två män i orangea overaller går längs en gata.
En man sitter med ett papper i sina händer.
Den stora bruna hunden hoppar in i en pool.
Tre personer står i en kylig juicegång i en affär.
En ung flicka lägger en liten bild i ett skumbakverk.
Lilla flicka med blå ögon äter kakor.
Fem personer hoppar i luften för en fotomöjlighet framför en fontän.
En grupp unga män delar ut i en park med sina skateboards.
En grupp människor äter på en restaurang med en väggmålning av en dam som handlar bakom sig.
En liten pojke, som är målad som en zombie klättrar på en stenstruktur.
2 kvinnor på en soffa, kvinna i vitt verkar beskriva något i hennes hand.
Border collie hoppar i luften och fångar en tennisboll.
En kvinna poserar med solglasögon formade som dollarskyltar och en silver resväska märkt "Lucky" full av sedlar.
En blond tjej uppträder karate och sparkar genom block av trä.
En person som bär hård hatt cyklar på gatan.
En halv naken man som hoppar ner i en vattensamling.
En byggnadsarbetare som pekar på ett föremål eller område som inte syns på bilden.
En liten flicka rider på framsidan av en kundvagn i en butik.
En kvinna i blå och vit skjorta bär cowboyhatt.
Kvinna med mörka glasögon och bollmössa som pratar på en mobiltelefon
Fågelns syn på en stadsarbetare som går på gatan.
Man rider JAL-bilen på en flygplats.
En ung pojke leker i en gul tunnel på en lekplats.
En kvinna med långt blont hår sträcker sig in i baksätet på sin bil.
En blondhårig pojke i röd skjorta och blå shorts som målar på en duk.
En pojke glider ner för en uppblåsbar vattenrutschbana.
Flickan i klänning hoppar i luften utanför.
Två kvinnor konsulterar en inköpslista medan de stannar i slutet av en gång på Target.
En liten pojke som sitter ute på uteplatsen och målar en bild.
En kvinna som går genom en parkeringsplats utan skor.
En äldre kvinna sitter nära en liten julgran med en olindad present och bär en lampskärm på huvudet.
Trädgårdsarbete är roligt och avkopplande.
Två kvinnor kickboxar, kvinnan i rött blockerar en kick från den andra leende kvinnan i blått.
En hund tappar en röd skiva på en strand.
Fyra tonåringar har en explosion i en källare spelar TV-spelet Rock Band.
En kvinna i röd skjorta med en mobiltelefon.
Två tjejer i en publik är klädda upp, en som den tecknade karaktären Wall-E.
Folk samtalar vid ett matbord under ett tak.
En brud och brudgum, klädda i leis, skär sin bröllopstårta.
Manliga hejaklacksledare håller upp kvinnliga hejaklacksledare på en fotbollsplan.
En grupp män som bär färggranna kläder twirl batonger unisont.
En liten pojke spillde sin mjölk från den gröna koppen.
En man står på toppen av en stenig kulle.
En mörkhårig man sköter en fruktaffär.
En kille med svart skjorta som sitter vid bordet och jobbar med datorprojekt.
String orkester och dirigent i rampljuset omgiven av mörker.
En man grillar korv medan två andra män äter i bakgrunden.
En mor och hennes sol sitter utanför.
En kvinna håller ett barn medan han läser.
Två män pratar medan de sitter på uteplatsen.
En grupp människor som sitter vid ett utomhusbord och äter mat och dricker alkoholhaltiga drycker.
Pojken med skjortan ogjord sträcker armen i luften.
En ung pojke i randig skjorta lutar sig mot ett träd medan ett annat barn sitter vid ett picknickbord.
Stranden med en person i en röd tanktopp som sitter under ett litet träd.
En rödskjortad man renoverar sitt kök, förbereder väggen bakom där hans disk ska sitta.
En pojke hoppar på en uppblåsbar vattenrutschbana
En man kastas av en häst på en rodeo.
En ung pojke som leker i en simbassäng
En äldre pojke och en medelålders pojke som skrattar åt en datorskärm.
Ett barn stoppar smuts i munnen på honom.
Sex kvinnor väntar på att få använda en port-o-john på ett fält.
En man förbereder en drake för flygning.
Två kvinnor i tutu ́s och benvärmare stannar för en pratstund.
Barn leker språnggroda bredvid fontänen.
En ung flicka i rosa skjorta sträcker sig för att röra vid en grön ballong.
Kvinnan leder sin lilla hund genom en hinderbana.
Vi gillar denna trädgård och vi njuter varje kväll på sommaren.
En man med ryggsäck pratar med en kvinna i svart skjorta.
En kvinna shoppar efter en spistopp i en förbättringsbutik och har hittat en som hon tycker om.
En kvinna i lila topp och vit mössa som joggar längs vägen.
En rödhårig liten flicka i lila fiskar på en båt ute på en sjö.
En man går på en låg lina under ett träd.
En pojke sitter på en beige stol bredvid en uppstoppad SvampBob Squarepants.
En man som cyklade på piren.
En brun och vit greyhound med en röd nummer fem fångas i luften racing.
En kvinna som passerar stranden.
En grupp barn i en kyrkkällare leker maracas och tamburiner.
En svart hund springer runt en utomhuspool.
En leende person som bär en svart ärmlös skjorta slår en spik i ett trästycke.
En staty av en ängel monterad på sidan av en byggnad.
En liten flicka och pojke sitter på en trälåda och läser böcker.
En leende man i förarsätet i en bil vänder sig mot baksätet.
En pojke ler och simmar i blått vatten.
En röd bil är fast i en explosion.
En man går fram till ett konferensrum.
Personen hänger glidande vid solnedgången.
En flygande maskin med gult segel landar med industribyggnader i bakgrunden.
Folk på en fullsatt stadsgata.
Alla på gatan i stan verkar vara upptagna med att göra sin egen grej.
Ett barn och hennes mamma leker boll i en park.
En man i kamelfärgad jacka som står och tittar på stengången.
En man i ventilationsmask snider en riddare på en tegelvägg.
Tre män ser ut som två andra män skära upp en nygrillad gris i trädgården.
En man som fångar en fisk från en båt.
En grupp människor som står och sitter runt vad som ser ut som ett stadshus möte.
En grupp människor som sitter vid ett bord och äter och pratar.
En kvinna med spaghettistrappad skjorta och en skjortlös pojke med röda shorts leker med en stor checkerbräda.
Ett barn som äter en hämtmatslåda
En man tittar på medan ett barn spelar ett spel.
En kvinna som bär klänning går över gatan.
En äldre man i vit skjorta går ut ur en byggnad genom ett par trädörrar.
Två barn håller ballonger och en kvinna är på en trottoar med en bil till sidan.
Ett skjortlöst barn spelar på en "häst" gunga gjord av gummi medan han håller en kvinnas hand.
Tre barn njuter av lunch på en picknickbänk tillsammans.
En pojke med röd skjorta skjuter fyrverkerier från en vågvägg i vattnet.
En man böjer sig ner för att tända ett fyrverkeri nära en sjö.
Två äldre pojkar i huvtröja låg på en madrass i en affär när två yngre flickor tittar på.
En brun hund som springer över gräset.
En man står i sin lilla båt mitt i sjön.
Ett barn i lila gör ett skateboardtrick.
En grupp damer ska ha fest.
En kvinna pekar medan andra tar bilder.
En grå hund med blå ögon som ligger på en ljusblå matta och tuggar på något.
En stadsarbetare förbereder sig för att hugga ner ett träd.
En grupp vänner sätter sig ner för något att äta.
En pojke som leker utomhus på en glid och rutschkana.
En ung flicka i röd skjorta som träffar en tennisboll med rosa racket
En man som sitter på en bänk och tar en paus från bygget.
Ett stort vitt rör sänks på en släpvagn, medan två arbetare står och väntar.
En ung flicka håller ett gråtande spädbarn.
Tonåringen övar med svärd i ett gym med sitt lag.
En liten hund sitter på en persons böjda ben.
En präst som bär en liten blå väska går nerför gatan och pratar på en mobiltelefon.
En man häller en drink i ett glas, medan en kvinna tittar.
Pojken som går bär grå shorts och ingen skjorta.
En stor grupp människor hänger på en stor gräsmatta.
En man i en grå t-shirt skyfflar cement från en skottkärra.
En man i hatt gräver nära ett stängsel.
En man skär trä för att lägga till stängslet han är i mitten av byggnaden.
En man i cowboyhatt trampas på av en brun häst
En man i randig skjorta dansar framför ett band.
Ett barn som bär en blå bandanna leker med en uppsättning färgade ringar.
Två personer forsar nerför en flod, en gångbro i bakgrunden.
Två personer i en kanot flyter förbi en stenig, skogbevuxen klippa.
En kvinna med blå blus och blå jeans rider i en cykel
Nån i grön skjorta som springer bakom en liten hund.
Kvinnan bär en lila skjorta och springer på stranden.
Ett äldre par sitter utanför en restaurang och njuter av vin.
En man i röd skjorta och en man i gul skjorta hukar sig i en skara människor.
En man som hamrar in en spik i en bjälke.
Två bruna hundar jagar och leker med varandra på sandstranden.
En dam korthårig dam med en tom tank topp tar bilder.
En grupp barn utanför en byggnad inkluderar en pojke som hoppar i gräset.
Två män under paraplyer på en gårdsförsäljning.
En man flyter på en liten båt nerför en vattengata i staden.
Kvinnan på stranden med en liten flicka.
Två gamla män med hattar står mellan bilar med dragspel.
En ung pojke tar bort ansiktet från en blåbärspaj.
En pojke sparkar en jättebaseball medan en grupp barn tittar.
En valp håller på att torka med en torktumlare
Ett litet barn i en rosa huvtröja stiger höga trappor utomhus.
En liten pojke hoppar ur poolen.
En söt brunett flicka lutar sig med handen mot väggen.
Två unga kvinnor står vid en Red Bull bil.
En kvinna som bär en bunt på huvudet leder två åsnor på en lerig gata.
Pappa njuter med sin i poolen.
En kvinna som bär en blå rutig skjorta tar mat från en gryta.
En liten hund som jagar en boll.
En liten pojke äter en klubba och dansar på gatan.
En grönskjortad man sitter bland de många obebodda röda sätena.
En skjortlös man har ett samtal med en sittande man medan en blond kvinna sover.
En baseballskytt som håller ett slagträ på fall.
En grupp shoppare kantar gatan i ett kommersiellt distrikt vid ett berg.
En man som sitter vid ett bord med en yxa och tittar på en trasig mugg.
En man står på scen med sin gitarr.
En far knuffar sina döttrar gokart medan en annan flicka tittar
En dam med hatt sittande framför sitt hus teckna porträtt
En kampsportartist bryter is med en spark.
En man som låg på marken i gräset omgiven av träd.
Tre kvinnor väntar på flygplatsen med sitt bagage.
En hund springer bakom en annan i en park.
Ett barn i en affär håller ett par betar mot kinderna.
En leende kvinna spelar fiol framför en turkos bakgrund.
Fyra män sitter i ett rum och tittar på någon.
Folk i vita skjortor och ryggsäckar ser sig omkring i en av dem med en liten kamera.
Två kvinnor solbadar vid vattnet.
Blå krabbor säljs från en hink på en fiskmarknad.
En cowboy och hans häst faller båda till marken på en arena.
En man som försöker hålla ut, när han tävlar i en rodeo på hästryggen.
En ung pojke står vid en bil som tvättas.
En man ser marken när han kommer in för en landning från parasailing.
Man försöker leda ett kit i öknen.
En man som pratar med andra män bakom en kamera på ett stativ.
Man går på trottoaren medan man pratar i telefon.
En pojke i gul regnrock undersöker en bit mat han håller i handen.
En man med långt hår sitter på soffan.
En man i röda shorts träffar en volleyboll i luften när en annan man tittar på.
En man med ryggsäck som går längs en väg.
Folk på en trottoar tittar in i skyltfönster medan andra bara fortsätter att gå.
En flicka går på en sandig stig.
En grupp människor går framför en tunnelbanebana.
En grupp människor som sitter utomhus.
En flicka i rosa byxor som springer, en utsmyckad spansk ruin i bakgrunden.
En tonåring i röd skjorta förbereder sig för att servera en volleyboll.
En kvinna står med ett barn bredvid en staty.
En brun hund som ammar
En lekfull hund hoppar på sanden.
En kvinna i röd skjorta med upplyft arm.
Tjej i blå tröja och håller en multicolor leksak sitter på axlarna på en man med grått hår.
En man i gammal kostym hoppar över en engelsk gata förutom en Peugeot.
Det finns tre män som bär kläder och står runt.
Två personer sitter på en bänk medan andra på avstånd rör sig.
En ung flicka i en röd plastbil i en fin skoaffär.
En man och kvinnor klättrar.
En ung asiatisk pojke i en orange långärmad t-shirt har en tidning.
En brudtärna i en knälång blå klänning går nerför gången med en brudgumman.
En man i gul slips och skjorta gör "hook'em horn" skylten.
En kvinna och en man står tillsammans.
En brud och brudgummen dansar i bröllopsmottagningen.
Brud äter bröllopstårta från sin nye mans skjorta.
En blond kvinna som bär en blå och rosa blommig bikini på en strand, redo att sätta en flaggstång i sanden.
Fyra män och en ung pojke sitter vid ett bord för trähantverk.
Ett barn kryper på ett trägolv nära en flaska vatten.
En liten pojke i blått kryper längs en fönsterbräda.
En man hjälper en ung pojke i en hatt att bygga något av trä med en hammare.
Ett barn i en ullmössa tittar på en låda.
En man som är utrustad med motorsåg och skyddsutrustning gör en fågelstaty av trä.
Två flickor ombord på en nöjespark.
En mycket attraktiv kvinna poserar framför en vacker växt under en solig dag.
Ett äldre par står i ett kök tillsammans.
Fyra personer står bakom en balkong framför en tegelbyggnad.
Ett blond barn inuti en låda som ler
En grön Volkswagen Bug och andra vintage bilar beundras av människor på en innergård.
Flera unga män surfar på C.D.
En grupp barn klättrar på en staty av en björn.
En äldre gentlemän sätter på sig ett enmansband med olika instrument.
En ung flicka sitter på skogsgolvet och tittar upp genom kikaren.
En kvinna rider en röd cykel längs en flod medan hon bär hjälm.
En infödd amerikansk kvinna som bär en färgglad skjorta arbetar på en vävstol.
En svart hund och en vit hund brottas.
En man klättrar över snötäckta klippor vid en strand.
En man som breakdansar på ett klinkergolv
Ett barn sover i en grön barnvagn.
Ett varuhus som säljer utländsk mat.
Många människor runt några lådor med fisk.
Tre bruna hundar springer efter en tennisboll.
En ung pojke ler när han hänger på apbarer.
Tre barn springer på gångvägen vid floden.
Den här kvinnan tar en paus efter en lång promenad eller joggingtur.
En grupp cyklister rider uppför gatan.
En svart hund springer parallell till ett stängsel i en gräsbevuxen medow.
En hund som springer med ett rött föremål i munnen.
Barn leker i det blå och gröna hopptältet fyllt med luft.
En man som jobbar under ett tåg.
En man med kamera med blå skjorta och jeans står mellan två höga byggnader.
Två pojkar leker i smutsigt vatten
En collegestudent messar ett meddelande till sin pojkvän medan hon väntar på att nästa lektion ska börja.
Äldre män gör sig redo för grillning.
En stor tunn hund springer snabbt i ett gräsfält.
En grupp män som bär röda och gula promenader.
En ung pojke sitter vid ett bord och äter som mat spills runt omkring.
Två arbetare i neongröna skjortor som öppnar en brukslåda.
En tonårstjej bär brun hatt och en jacka med hjärtan på.
Den här unga flickan njuter av barndomens oskuld och det varma vädret.
En ung kvinna, klädd i avslappnat svarta kläder, håller i ett svärd, i stridsställning.
Barn i sommarkläder spelar på en turnaround i en soldränkt park.
Greyhounds springer snabbt i det här loppet.
En grupp människor går omkring utomhus, en flicka bärs.
Denna kyrkokör sjunger för massorna när de sjunger glada sånger ur boken i en kyrka.
En man står bredvid ett tåg.
2 unga flickor sitter framför en bokhylla och 1 läser en bok.
Ungar hoppar från en pire i vattnet i skymningen.
Ett par på vägkanten som pratar.
En liten vit och brun hund hoppar över en horisontell stolpe.
En brun och vit hund som simmar mot några i poolen
En man i vit skjorta som gräver ett hål.
Barn sitter vid ett långt blått bord och ritar bilder med kritor.
En äldre person och ett litet barn går tillsammans framför en stor byggnad.
En kvinna i blå topp och hatt sträcker eller utför yoga på stranden.
En man som bär skyddskläder slipar ner ett stort metallföremål.
En svart hund i ett plant fält försöker göra en sväng.
Pojkar i uniform bakom en boll.
En kvinna med grön topp åker rullskridskor genom en folkmassa.
En man sitter på en cykel fäst vid en pelare i luften.
En ung man i udda kläder lutar sig mot en tegelvägg med en trädgård i.
En ung flicka njuter av en frusen behandling vid poolen.
En fotograf knäböjer bredvid kanten av en docka med sin kamera.
Två män tittar mot marken medan en bär handskar och håller i ett verktyg.
En ung man spelar elcello framför en kvinna.
En man som bär glasögon spelar gitarr framför en mikrofon.
En man i badbyxor kramar en kvinna i cutoffs och en bikini övredel i en fontän.
En man med bröd som tittar på kameran.
Två hundar, en kommer mot kameran medan en går i bakgrunden.
Den lilla flickan har en lila klänning på sig.
Flera kvinnor i huvudskarvar står på en kullerstensgård.
En flicka och en pojke sitter på marken omgiven av växter.
Den svarta och bruna hunden står med benen isär på stranden.
En man med en kopp framför en träkonstruktion.
En ung topless man som bär solglasögon och shorts håller i en fotboll.
En liten hund hoppar några hinder.
Två män, två barn och en kvinna som alla sitter nära en monter fylld med väskor.
Tre män går tillsammans på en plaza.
En ung man med shorts och ingen skjorta är hög sparkar som vatten flyger från hans kläder.
Fem stråkmusiker spelar tillsammans på en scen.
Tre män i svarta kostymer tittar på något framför dem.
En äldre kvinna med käpp i solglasögon sitter på en bänk.
En äldre asiatisk man i blå rock med käpp sitter utanför en tegel- och cementbyggnad äldre.
Folk som sitter utanför under ett grönt paraply.
En svart hund, i en Alley kanske, Han kan vara vilse, och Cold, eller Hungry.
Man och kvinna som bär svart gå med armar runt varandra.
En ung flicka sitter på trottoaren och byter däck på en cykel medan en annan ung flicka sitter och tittar på henne.
Ett barn ligger i en sandlåda och leker med en hink.
Den unga damen verkar vara en mimare bland sina kamrater.
En fet kille i rosa som dricker öl.
En hona i blå jeansshorts och en svart topp som sitter i en korgstol.
En liten hund hoppar över ett hopp.
Äldre man som spelar ett udda gitarrliknande instrument i vad som verkar vara en park eller ett öppet område.
Ett barn leker i vatten på gatan.
Tre män är på väg in i en byggnad på väg tillbaka till arbetet.
Flickan utanför håller en rosa blomma som matchar hennes topp och leende.
Flera personer förbereder sina stånd som består av fisk, grönsaker och frukt för det allmänna ögat.
En man med blå skjorta och hatt hoppar på ett hjul på en fontän avsats
En man går genom en byggnad och håller ett litet barns hand.
Den store mannen tar en plats på en restaurang.
Fyra personer, tre flickor, en pojke, sitter i en båt.
En hona med glasögon, en brun skjorta och en ryggsäck.
Elva personer står på en balkong och tittar ut över träden och faunan utanför.
Ett europeiskt par som står på gatan och kysser varandra.
Hund och kvinnor med barnvagn korsar en bro på landsbygden.
Man leker hämta med sin hund nära en båt docka.
Två små vita hundar leker ute i snön.
En skara kvinnor är inblandade i en opinionsbildande promenad.
Två barn sitter i en barnvagn framför en brandbil.
Två män i hattar spelar banjo och saxofon utomhus med en hattad man som sitter på en bänk bakom.
Ett litet barn med grå skjorta och napp står bredvid en leksakshäst.
En kvinna i svart skjorta går nerför gatan
En vit hund med svarta fläckar springer genom en spray från en slang till en blå plast vaddbassäng.
Akrobatiska underhållare utan skjortor uppträder för åskådare.
En tonåring hoppar högt på en studsmatta och ett litet barn faller på hans mage.
En grupp människor tittar på en flerfärgad bild på en skärm.
Kvinnan med en hennatatuering håller ett papper i sin vänstra hand.
En grupp människor gör sig av med en berg-och dalbana.
En kille i blå skjorta bredvid en man i vit skjorta som tittar på en kille i orange skjorta.
Kvinnan står och tittar på rader av tidskrifter.
En asiatisk kvinna som bär en blå rock och rosa tröja håller upp en silverpärla för att undersöka den.
En massa människor går nerför en trappa.
Flera personer pratar och dricker öl medan de sitter vid ett picknickbord.
En äldre asiatisk man, klädd i orange rock i storstadsområdet.
En man med ett ansikte målat som en clown bär en cowboyhatt.
Flickan snurrar långa, färgstarka streamers.
En äldre man som reparerar en skrivmaskin omgiven av andra skrivmaskiner.
Små flickor sover på golvet.
Höger ben i en tandställning, en ung pojke ligger på soffan medan han använder sin mobiltelefon.
Folk sitter och klättrar på stora klippformationer.
Tre blonda tjejer och en mörkhårig tjej försöker sälja dekorerade skal och stenar.
Två personer tillagar en måltid tillsammans i ett kök.
En liten pojke som bär en brun t-shirt suger på en nappare med handen i luften.
Fyra unga pojkar som böjer sig för kameran.
En ung asiatisk kvinna i orange klänning som pratar med någon.
En häst tjänar pengar på sin ryttare på en arena som åskådare tittar på från blekare.
En indisk man står bland en grupp indianer som skriver på en skrivtavla.
Lilla flicka bär massor av rosa leker med sin cykel.
Få barn cyklar runt en stig med shorts.
En vit hund som kommer ut ur en blå tunnel.
En man i vita byxor som går genom en arbour av människor som är vända mot varandra sammankopplade med sina händer.
En man klädd i orange ser ut som han spelar ett instrument.
En brun och svart hund som ligger bredvid en färgglad boll.
En pojke leker med en nudel vid poolen.
Två små barn som har kul på en berg-och dalbana
En kvinna är svart och valvar.
Två kvinnor i röda kjolar som dansar för en publik.
Man och två barn på en båt på sjön.
En grupp människor sitter på stranden, bortom ett tecken som varnar för oseriösa vågor.
Två små flickor som svänger sida vid sida i en park på en varm dag.
En grupp människor sitter under en parasoll i en gräsbevuxen skogsglänta.
Två honor i kjol går på trottoaren.
En blond kvinna i grissvans går nerför trottoaren barfota med en grön tub på ryggen.
Kvinnan hukar sig mot en tegelvägg och pratar på sin mobil.
En man i solglasögon skriver på en pad med sin cykel lutad mot honom.
Mannen har en svart och vit halsduk runt halsen.
En kvinna i röd skjorta och en man i vitt står framför en spegel.
En grupp barn i tonåren går nära en flod.
En man med mustasch håller två pojkar i en pool.
Närbild av person som spelar en marsch band snara trummor.
En hund uppträder på en hundutställning.
Unga pojkar som spelar Wii.
En baseballspelare i uniform som precis kastade en boll.
Två personer på en surfbräda i vattnet
Lilla blonda flicka som kliver på en blå yta utanför.
4 personer går genom öknen.
En brun hund springer över gräset med en käpp i munnen.
En hund jagar en fågel i vattnet.
Människor åker skridskor i en urban utomhus skridskobana
En man åker skridskor på en järnväg.
En man utan skjorta poserar med armarna utspridda bredvid en kvinna.
En liten pojke som bär pyjamas vänder äggplantan på gasgrillen.
En grupp vuxna leds av en äldre gentleman i en övning med gruppansträngning för att stabilisera en lång stav.
En ung man i GIGOLO-skjorta vid receptionen.
En ung flicka i röd baddräkt simmar i en pool.
Hunden rinner genom vattnet på en strand.
En flicka är vänd mot en vägg med ryggen mot ett kupolliknande konstverk.
Tre rugbyspelare försöker fånga bollen
De tre männen hoppade i luften i ett försök att ta bollen.
En lånelöpare deltar i ett lopp i regnet.
En kvinna i rosa skjorta som står framför en gul byggnad.
Två vuxna sitter på en bänk.
En person med en elektrisk borr som gör något mot ett leksaksdjur.
En man ler medan han håller i ett gråtande spädbarn.
Mannen med rakat huvud och piercingar i bröstvårtan bär solglasögon.
Ett barn springer nära några träd.
En brun och vit hund springer snabbt på en inhägnad gård.
Två flickor tittar genom ett mikroskop.
En svart och brun hund springer och plaskar i vattnet.
Fotboll spel med lag i rött och blått.
En man i vit skjorta glider genom sanden mot en man i blå uniform och hatt som håller ut en sporthandske mot honom.
Man med skägg gör skateboard stunt
Ett par spelar frisbee i ett grönt fält med träd i bakgrunden
En kvinna i en blå skjorta som sköljer ut sin mopp på gatan.
En man, klädd i en vit knapp ner skjorta och glasögon, skriver på en bärbar dator.
En äldre man lagar korv på en grill.
En vit kvinna och en svart man i en röd hatt spela slåss.
En flicka och en pojke begraver en annan pojke i sanden.
En kille med en rosa skjorta som sitter på marken och ritar en påfågel med krita.
Hundar i vattnet med en basketboll och en person på hästryggen.
Barnet sover i en spjälsäng med tändstickor, en elektrisk borr och några uppstoppade djur.
En svart hund biter på en fotbollsboll på marken.
En exalterad pojke som leker i surfingen med en kroppsbräda.
Pojken vadar genom det blå havet.
Ett barn med tandställning och en blå hatt visar botten av sin skateboard.
Det finns en chun kuk do turnering med en grupp åskådare tittar på.
Två kvinnor sparrar våldsamt på Tae Kwon Do konkurrens, medan domare klockor.
Ett band uppträder på scenen.
Det finns ett barn runt 6 månader gammal sitter på en stor Elmo docka, ser ut som han är på väg att tuggummi den med en Sesam Street bok i sin högra hand.
En beagle klättrar genom några grå trappor.
En man och en kvinna i baddräkt håller varandra i en vattensamling.
Deprimerad man som inte vet vad man ska göra.
En kvinna som bär en röd och vit klänning har en lång halsduk bakom sig.
Tre forskare som arbetar i ett labb.
Tre barn springer framför sin mamma i en park.
Tre barn åker skridskor på rullskridskor.
En brun och vit hund leker i en pool med en man.
En fårhund föder upp får på en gräsbevuxen stig.
Två hundar i en röd bil som tittar på en kvinna som kliver ur sin bil.
En flicka skakar upp vattnet ur håret.
Fyra unga män sitter på golvet nära en TV som visar Elmo från Sesam Street.
Äldre vuxna och unga vuxna, ha fest och dansa.
En grupp människor i en cirkel klappar händerna medan andra sitter i bakgrunden.
Tre unga män spelar domino medan en äldre kvinna tittar.
En man i blå skjorta och sandaler kastar ett föremål mot ett mål medan en grupp äldre vuxna ser på.
Amputerade stående från rullstol kasta en boll i en senior center.
En man i orange skjorta håller ett föremål och talar med en flicka i en blå skjorta som tittar tillbaka på honom.
Två män bestämmer vad de ska göra med en blockerande fallen gren.
En ung man i röd randig skjorta och blå jeans bowlar med en blå boll i en bowlinghall.
En grupp individer sitter i ett rum tillsammans och ler.
Män arbetar i viss vegetation bredvid en tegelstruktur.
En person spelar på apbarer medan andra tittar.
Två män står på taket av en hög betongkonstruktion.
En tonåring sitter väldigt högt i ett träd.
2 personer står upp klädd i svart på en gammal persons hem, medan några åskådare sitter i rullstolar i närheten.
Tonåringar interagerar med äldre människor i ett gemensamt rum.
En gammal man dansar bara med en kvinna.
Två flickor, en i röd skjorta och blå kjol, tvättar en röd lastbil.
En grupp på 8 tonåringar som sitter längs en vägg och håller i ett snöre.
Två män deltar i en blandad kampsport tävling.
En ung kvinna som bär en rosa och grön randig skjorta med ett vitt bälte och flip-flops sittande på ett cementsteg.
En svart hund med blå krage går genom det gröna gräset.
Tre barn står runt en figur på ett lila bord, två barn har vita rockar på.
En kille som spelar basket med åskådare som tittar.
En man i svart mössa tittar bort från en kvinna i svart och vit polka-prickad klädsel.
En man i svart skjorta som dansar med en kvinna som ler.
Två män byter korv med varandra via munnen.
En man gnager efter äpplen i en plasthink.
En grupp tonåringar sitter i en cirkel; mannen i mitten sitter på golvet och det finns en kvast som står bakom honom.
En kvinna organiserar sin mat i mjölkkorgar.
En kvinna har många kartonger med olika livsmedel utanför och håller en burk.
En ung man i jeans och en röd skjorta, klädd i gula handskar, håller i en trädgren.
Tre personer står högst upp i en utomhustrappa.
En kvinna tittar som sin vän går för en reserv.
En man som håller i en kofot och bär masker ser upp.
Två flickor hjälper till att städa ett smutsigt hus
Tre personer städar fönster och en kvinna i en blå skjorta pratar med dem.
En man filmar en grupp flickor utomhus.
En fisheye lins fångar en ung flicka med mörkt hår på lekplatsen.
En äldre kvinna och en ung man spelar bingo.
En kvinna har en "biltvätt" skylt på kanten av en lugn gata.
En man i brun skjorta och blå shorts som går i Droney Park.
Några pojkar och flickor sitter ner i en nöjespark rida.
Tre barn leker i en yttre träkonstruktion.
Några män sitter utanför ett område med en öppen grind äter sina luncher.
Flera barn tittar på karneval spel.
Två flickor i denim shorts står i en pöl med vatten.
Två unga barn springer på sand mot en stor vattensamling.
Två hanar och en hona som leker i en källa med vatten.
Ett barn och golv täckt med vitt pulver.
Två personer med djurtryckta byxor som ligger på en säng bredvid varandra.
En hund springer genom högt gräs.
Hunden springer i gräset med en leksak i munnen
Två tävlande cyklister trampar förbi åskådarskaror.
En man sitter framför en vägg med konstbilder på sig.
Två rödhåriga pojkar med glasögon står på bänken och slåss med pinnar.
En flicka i en färgstark hatt har en konstig varelse som vilar på hennes hand.
En liten grå hund hoppar över ett litet hinder.
En man står på toppen av en glaciär.
En ryttare på en häst framför en bergskedja
En grupp människor i ett cykellopp.
En man i rosa skjorta rider en häst.
En tjurryttare rider en tjur medan andra cowboys tittar på och väntar på att hjälpa honom om det behövs.
Ett barn glider ner för en grön rutschkana.
Kid i Jean shorts använder en skateboard för att hoppa över en kameraman medan andra skateboardare och kameramän klockor.
Två långa svarta hundar springer genom högt gräs.
Kvinnan bär en svart hatt med en amerikansk flagga på.
En kvinna som går in i vågorna.
En person i shorts håller en Frisbee medan teammedlem i röda skjortor och åskådare tittar på.
En ung vuxen i svart skjorta sticker handen i en djurfälla.
En man på en arena som försöker stanna på en häst så länge han kan.
En man med mohawk ler mot kameran.
Flera hundar springer ut, med två fordon i bakgrunden.
Tre skällande, ylande hundar
En brun hund i luften med en frisbee i munnen.
En man som sprutar en superdämpare i munnen på en hund.
Barefoot människor står i vatten framför ett stort konstverk med ett ansikte.
En kvinna som balanserar ett svärd på huvudet.
En svart och vit hund hoppar genom luften när två människor tittar i bakgrunden.
En man i en coca cola byggnad torkar ner ett bord.
En tjej basketspelare klädd i blått blockerar en annan tjejspelare klädd i gult.
Människan står på kanten av klippor nära ett hav.
Två personer dyker i det blå havet.
Två pojkar tittar genom ett fönster på en flygplats.
Två små barn leker i en barnpool med vattenkanoner.
En stor, ståtlig stadsstaty på natten.
Kvinnan stänker vatten ur en hink.
En man i blå skjorta och vit hatt som städar en fontän.
En man med svart rock och röd hatt håller en kamera.
En man i vit skjorta kysser en liten pojke när han håller honom.
En stor skåpbil kör ner för en nationell väg i höst.
Ett marschband i full uniform kommer nerför gatan.
En unge i vit skjorta är i ett högt träd.
En liten flicka som håller i en glasstrut och slickar på läpparna.
En kvinna sveper sina armar runt en man när han lutar sig in för att kyssa henne.
En man i vadare fiskar efter något i en pool.
En kvinna har två barn att ta hand om medan hon är ute, en sitter på axlarna och den andra sitter i hennes knä.
En blond kvinna i svarta jeans sitter på en vägg och undersöker naglarna.
Kvinnan håller i en mugg och har solglasögon på huvudet.
En man som tar en tupplur på en varm eftermiddag.
På havssidan joggar en flicka i gula byxor och en pojke som cyklar.
Fyra barn leker runt en stolpe.
En svart och vit hund som leker med en vit boll i ett glest brunt fält.
En vit hund springer på stranden.
Två hundar leker och brottas med varandra.
Ung pojke med glasögon som leker i sprinklern.
En grupp kvinnor går nerför en gata på natten.
En man tittar på en skulptur i ett stort tomt rum.
En man med rakat huvud och solglasögon ler brett.
En tjej i vit klänning och röd väska som pratar i telefon.
En ung flicka och en ung man som spelar kastspel på en utomhusfest.
En rödhårig pojke med glasögon som blåser i en stor bubbla
Ung man med en svart skjorta på, rider en blå cykel med en baby som sitter framför honom.
En man balanserar en tallrik mat på huvudet.
En kock lagar mat medan två tittar på.
Folk står på båtbryggan och väntar på att deras båt ska komma.
En man som bär en orange väska går förbi två telefonlådor i brittisk stil.
Två barn slåss på ett torg medan folk tittar på.
En publik samlas för att se två män uppträda en brasiliansk dans.
Flera barn står framför en byggnad.
En varierad grupp individer sitter på en gräsmatta på sommaren.
En skjortlös man åker på sin skateboard medan han går sin hund.
En lurvig hund hoppar över ett hinder.
En pojke med mohawk och solglasögon.
En man och kvinna som bär solglasögon och vita t-shirts ler för kameran.
En ung pojke tar ett bad från en hink.
En man med långt hår bakbunden och bär en blå skjorta spelar klarinett.
En skjortlös man som sitter på en sten vid en blå byggnad.
De två pojkarna leker ute på fältet.
Två personer ligger i en säng mitt i ett varuhus.
Två personer, med byggnader bakom sig, står nära en blå bil med två dörrar öppna.
En tysk korthårig pekare vilar på en matta vid ett soligt fönster.
Två stora, svarta hundar leker med en kollapsad boll.
En liten pojke hoppar in i barnpoolen i trädgården.
Ett barn i baddräkt leker i en sprinkler.
En vit hund springer mot kameran när en man går sin väg.
Arbetare som drar ett rep fastsatt i vad som verkar vara en båt.
En dam med blont hår som hjälper en annan person.
Tre mörkhåriga människor står nära varandra med stora byggnader i bakgrunden.
Jag ska till en korvtävling på Coney Island.
En grupp tjurar springer längs en gata när folk springer och andra tittar.
En tjej som bär solglasögon ler för kameran.
En kille som gör tricks på en motorcykel.
En motorcykelförare står ovanpå sin cykel.
En ung pojke ligger i vattnet vid stranden.
Två tonåringar på stranden leker i sanden
En ung asiatisk man och kvinna som satt framför trappan på ett litet företag och rökte cigaretter.
Två unga pojkar leker med ett pussel i ett klassrum.
En fotbollsspelare fick ett pass medan de två spelarna från det motsatta laget försöker märka honom medan han är på marken.
En grupp kaukasiska människor som ligger i ett sandigt område.
En ung man hoppar ner i vattnet från en flytande rutschkana.
Två kvinnor som plockar växter i en öppen dal.
En svart hund med ett band på står framför några andra prisband.
En man som fotograferar med hjälp av sina zoomlinser.
En liten flicka med hästsvans skrattar nära en plast slott spela uppsättning.
Ryttaren kastar upp handen för balans som de bruna hästpengarna.
En kille i en Nike-skjorta som läser "MAKA NÅGOT BULLER" lutar huvudet i sidled när han äter.
En man i korta shorts poserar på en stor sten.
Den här kvinnan bär en vit t-shirt och håller i en kopp.
En grupp män går mellan järnvägsspåren.
En grupp klädda upp människor tittar på en broschyr försöker bestämma vilken webbplats att se nästa.
En man med bandage på fingret klättrar som andra tittar på.
En grupp barn sitter på golvet mot en tegelvägg medan en kvinna iakttar dem.
En äldre man som sitter vid en upplyst arbetsbänk.
En leende kvinna i bikini i luften över en dykbräda.
En man förbereder sig för att slå en backhand tennis shot.
Två små pojkar med målade ansikten sitter bredvid varandra.
En grupp tjejer på en strand.
Två unga flickor, en blondin och den andra brunetten, hoppar på en grön soffa i ett ljust, soldränkt rum.
En man i röd skjorta spelar tennis utomhus.
Man i mitten steg upphängd i luften, på väg att svinga en tennisracket på en tennisbana.
En musiker på trottoarkanten som visar sin talang offentligt.
En man i blå skjorta läser ett papper.
En man i förkläde ler när han pommes frites mat.
Två kvinnor sitter vid några stenar medan en av dem dricker.
En kvinna som går med ett blått paraply.
En ung man står på en rulltrappa med en kamera i handen och tittar blankt in i bilden.
En leende liten pojke hoppar upp till en leksak basketkorg.
Två unga flickor i klänningar står tillsammans framför en gul vägg.
En baseballspelare som träffar en boll.
En brun hund och en svart hund leker med en leksak.
Den här flickan plockar blomman från växten.
En grupp människor står längst fram i rummet och förbereder sig för att sjunga.
Några killar som dansar en ceremoniell dans i en parad
En mycket glad baby i en gul skjorta som svänger på gungan.
En kvinna med en speciell typ av cykel tittar på ett barn.
En tjej i bikini som börjar få slut på surfing.
Kvinnan i tanktoppen har en tatuering på armen.
Mike Holmgren på fältet med sitt lag Seattle Seahawkss pratar om övningsdetaljer med en assisterande tränare.
Folk hoppar från en mycket hög bro ner i vattnet nedanför.
En äldre man höjer sitt vinglas under en utomhusmåltid med andra.
En kvinna i röd klänning tittar ut genom ett fönster.
Två små pojkar spelar ett spel, en med munnen vidöppen.
En tränare som bär en blå skjorta pekar ut en kamera.
En man i hundkläder spelar vid ett kortbord med en illasinnad kvinna och langare.
En liten pojke jagar duvor på gatan och en man tittar på honom.
En man och en kvinna ses kyssas nära ett öppet fönster.
En grupp kvinnor kramar varandra
En vit hund som får godis i munnen.
En man som sitter på ett räcke på en konsert.
Många människor samlas i olika delar av en gammal byggnad.
En mogen kvinna i solglasögon och en jeansjacka.
En man paddlar en båt medan fyra kvinnor står på en sten i en vattenförekomst
En pojke hänger upp och ner från en metallstång.
En svart och en brun hund som springer i gräset.
Två pojkar leker med två hundar på stranden.
En ung kvinna med en blå Mohawk ser åt höger medan hon håller i en liten hand som tittar åt vänster.
En ung flicka i baddräkt som åker leksakståg.
Fyra flickor lagar mat på ett bord utomhus.
En man hoppar framför ett palats i Kina.
En svart och vit hund springer i gräset.
En man tittar i fjärran bredvid en annan som har sin hand i luften.
Modern med två söner simmar i havet.
Fem barn sitter på en trätrappa och poserar för en bild.
I skogen förbereder sig en ung man med röda shorts för att kasta en frisbee.
Två fotbollsspelare stöter på varandra.
En flicka i rosa solklänning cyklar bredvid ett vitt staket.
Tre poliser samtalar med rullskridskor.
2 Manliga Camp Rådgivare koppla av under eftermiddagen ledig tid för sin ungdom som direktören talar om de kommande kvällsaktiviteter
Ett blond barn ligger på en gren av ett träd på ett grönt fält.
En kvinna i en sari bredvid en pojke som håller ett rött paraply på en regnig gata
Två män använder keramiska plattor på ett gammalt tak.
En hund står på bakbenen i ett skogsområde medan en annan hund tittar.
Den svarta hunden bär en limegrön krage.
Tre män i västar som sitter i närheten av en hög med smuts med ryggen vänd mot en vägg.
Den unge mannen väntar med andra på trottoaren.
En ung tonårspojke röker en cigarett framför ett järnstängsel.
Folk pratar på en asiatisk marknad.
Ett barn med en vattenpistol som sprutas med vatten.
Fyra artister är på scen och interagerar med publiken.
En blond tjej sitter och dricker läsk och tittar på en delfin som simmar i bakgrunden.
En kvinna i röd skjorta sjunger.
En man som går längs en gångväg i ett gäng butikslokaler.
Två stora hundar springer i lite gräs.
En man i en mössa putsar en växt utomhus.
En långhårig man framför mikrofoner med musikinstrument.
En man med slickat bakhår och svart rock spelar en bandspelare.
En ung kvinna målar ett skyddsräcke.
En grupp människor poserar för en bild av ett metallskyddsräcke.
En man som planterar blommor runt en stolpe utanför.
En man och kvinna gräver upp jord och har en växt nära dem.
Folk som sitter i stolar med en rad flaggor hängande över dem.
Antalet små barn är betydligt fler än de vuxna i matsalen.
Kvinna inför gardinerade fönster och glas renare samtidigt hålla en pappershandduk.
Kvinnan i en blå klänning med ett lila paraply stående på vägen.
En baseballspelare glider mot en bas.
En ung flicka sitter framför en utställning på ett akvarium när en delfin simmar förbi.
En kvinna står på trottoarkanten bredvid en livlig gata.
En man använder en proffssåg för att fixa gatan.
En publik tittar på en utomhuskonsert.
En kvinna som går framför en lastbil och pratar med någon som går bredvid henne.
Tre unga människor planterar blommor och täcker området med en presenning.
Människor planterar blommor utanför i en cirkel.
Två personer i röda skjortor städar en gränd.
En kvinna ler åt ett barn medan ett äldre par ser på.
Små barn skjuter korgar på fältet.
En man som sitter i en grön stol framför ett stort fönster och tittar ut mot en stadsbild.
Folk är på en restaurang och äter.
Solen skiner ljust på snön som omger några få människor.
En ung man bär brun hatt och solglasögon.
Kvinnan i röd skjorta och snygg tittar på småsaker vid ett bord.
En publik tittar på ett band som uppträder på trottoaren.
Fyra personer i ljusblått vatten med ett barn i en rosa inter tub.
Flera personer slutade vänta på att tåget skulle passera.
En grupp greyhoundhundar springer runt ett grusspår.
En pojke i gul skjorta som springer förbi några fåglar.
En man drar en massa smuts i en smal gränd där en motorcykel står parkerad.
Ett märkligt barn som försökte fiska vad naturen spolade i land med en vacker havsbakgrund.
En man som kör en orange och vit motorcykel.
Den blonda kvinnan håller i ett svart paraply.
En kvinna med käpp som bär påsen går längs trottoaren.
En ung indianmamma är med sitt barn.
En grupp arbetare på en strandpromenad bär fluorescerande västar och håller lätta trollstavar.
En grupp människor gör sig redo för att bestiga ett berg.
En liten hund leker med en plastpåse på trottoaren.
En liten hund hoppar över en gul bjälke.
En man som håller upp en liten flicka i luften utanför.
Folk använder datorterminalerna på ett modernt bibliotek.
3 män spelar och rider på ett fordon gjort av musikinstrument inklusive en trumma och ett piano.
En man valv över en hög bar.
En grupp ungdomar utgör en bild på ett område
En man i shorts spelar beachvolleyboll.
En ung flicka hoppas från sten till sten i sina bara fötter.
De här tjejerna har jätteroligt att leta efter snäckskal.
Två personer i ett tätt djungelområde med träd och gräs överallt.
Mannen i förklädet förbereder matbordet.
En liten pojke spanar en slang på sin bror som är på andra sidan fönstret.
Hundar tävlar runt en kurva i banan.
Flera förskolebarn står och tittar genom staketbarer när två vuxna tittar på.
En medelålders man skiner svarta läderskor.
En soffa sitter trasig medan en man sitter ett bord bakom dem.
En grupp människor står och lyssnar på en talare.
Ett barfota barn går på stranden mot havet.
Fyra hundar plaskar i vattnet
En man i randig skjorta poserar med en blond tjej i svart förkläde.
En hund som jagar en frisbee i vattnet
En kille som dricker ur en stor silvermugg, vars innehåll är okänt.
En liten flicka i rosa klänning går ut.
En asiatisk man som håller i ett stort antal väskor ser ut över en gata.
En kvinna med vit topp med design på framsidan som rengör det vita räcket.
En äldre man med händerna placerade på en tunna på en lastbilsgård.
En afrikansk amerikansk kvinna med två unga flickor.
Tre äldre män spelar livemusik i en stor sal.
Fyra tonåringar är i en kyrka och spelar sina instrument.
En man i senapsgul jacka sitter framför vattnet medan han läser.
Mannen spelar ett stränginstrument på marken.
Ett barn i en randig tank topp skateboards nerför gatan
En flicka i en skara som håller fast vid ett koppel får.
En man med cykelhjälm och två unga pojkar har bara huvudet kikat upp från en hög med löv.
Ett barn äter aqua-färgad tårta väldigt stökigt.
Två barn sitter utanför vid ett bord med popcorn över hela det.
En man med en blå jacka tittar på objekt.
En man med en vit krageskjorta på vattnet.
Ett par tar en paus från dansen.
En grupp människor, inklusive en barfota kvinna med vita shorts, en svart jacka och ryggsäck väntar på ett lätt tåg.
Två små pojkar leker i vattnet som sprinklern lämnat efter sig.
Två män sätter gips på en byggnad.
Ett barn leker i en mångfärgad fontän.
Ett barn flyter på en flotte och plaskar i en pool.
Man i vit jonglering med en cykel mot väggen.
Fyra pojkar kommer att drabbas av en annalkande våg.
En grupp människor står på trottoaren och tittar tvärs över gatan.
En man, klädd i vit t-shirt och jeans, sitter på två staplade lådor medan han spelar gitarr för tips.
En flicka svänger över vågorna på en repsving.
En liten flicka i gul skjorta springer genom en fontän i en livlig park
Ett band som spelar i en bar framför en publik.
Ett barn sitter på en rosa, blommande soffa och läser en bok.
Två kvinnor jobbar i ett kök.
Ett ungt barn med vilt lockigt hår sitter på en stol och visar upp sina legos.
En gatuartist och hans gitarr målade helt blå.
Två pojkar skateboardar framför en kontorsbyggnad.
Två män som spelar gitarr på scenen
En man störtar ner i vattnet med sin fallskärm.
En kvinna som hjälper ett barn ut ur poolen.
En kvinna, en pojke och en hund går uppför en kulle.
En man spelar golf och slår bollen ur en sandbunker.
En man i jeans sover med en röd mask som täcker hans ögon.
Det finns två greyhounds racing runt en grusspår.
En indisk hane dricker något ur en lerbägare.
Man tar en paus under ett paraply lutar mot lastbil.
En man i rosa skjorta och vita byxor i mitten av hoppet spelar gitarr.
Kvinnan på bänken tittar på molnig bergsutsikt.
Två kvinnor i sandaler, en i grön hatt binder den andra kvinnans klädband.
En kvinna i svart skjorta tittar på en cykel.
En kvinna i orange tröja håller ett glas i handen.
Två unga pojkar som dricker hemma.
Ett rockband spelar i en svagt upplyst bar.
En hund rullar i gräset.
En blondhårig pojke med röd skjorta och röda shorts som klättrar i ett träd.
En man står på en stege för att ta en bild med sin mobiltelefon.
Flera kvinnor som bär vita skor och sandaler går genom en gatufestival.
En man slår till ett städ.
En liten flicka erbjuder en boll till en upprörd småbarn på ett gräsrött fält medan en man i bermuda shorts står bakom dem.
Svart hund leker med en vit och blå leksak.
En man kör lastbil medan ett barn sitter i knät och styr.
Två unga flickor klädda i sin söndags bästa kamrat över ett staket.
En man går mot en polis som står på en trottoar på en stadsgata.
En man står på en trottoar mellan en gräs gräsmatta och byggnad
En man i vit skjorta och blå jeans som går över betong.
Kvinna som sorterar hink med mat.
En man ritar på gatan medan en annan man filmar det.
En man säljer mat på ett gatustånd.
Pojken sitter i bilens chaufförs knä och hjälper till att styra.
En kvinna visar en man något på sin mobil mitt på en fullsatt gata.
En grupp människor sitter bredvid varandra med en del vita skjortor och blå västar med gula stygn och de andra med stora fluffiga vita hattar med rosa fluffig topp.
Män och kvinnor i traditionella klänningar deltar något.
En liten pojke leker med en pistol på trottoaren utanför.
En kvinna jobbar på ett matställe i stan.
En person som hämtar något från en påse på en matlagningsdisk.
En gata med många annonser.
En asiatisk kvinna går till en pelare bredvid en byggnad.
En man gör sig redo att slå en tennisboll.
Ett barn i blå skjorta har ett armbandsur.
Två män sitter på motsatta sidor av en busshållplats
En man, kvinna och liten flicka går längs en strandpromenad vid ett lugnt hav.
En flintskallig man hjälper en ung pojkfisk.
Ett par njuter av utsikten över vattnet medan de sitter på en uteplats.
En man sitter i en stol medan han håller i en stor stolpe.
En grupp människor från Mellanöstern går genom snön.
En flicka som sitter på en mans knä på ett passagerartåg
Ett litet barn rör om i maten med en röd sked på köksdisken.
Hur tar vi oss till andra sidan?
Mannen och kvinnan kramar och kysser nära musiker som uppträder.
Den här kvinnan spelar ett instrument.
En hund hoppar över en buske på stranden.
En pojke hoppar från en hög klippa till vattnet nedanför.
En pojke går ombord i en bakgårdspool medan två andra vaktar.
En man som sjunger framför ett stort hjärta.
En hund hoppar för att försöka fånga en gul tennisboll på en uteplats.
En man böjer sig ner och gräver i en vit väska.
En kvinna som står framför en strandscen och ler.
En man med svarta glasögon spelar en svart gitarr.
Detta lilla barn sitter bakom ratten på en bil.
En hund springer iväg på sanden.
En ung flicka som visar sin lila tunga
En stor grupp människor samlades utanför.
Någon som står på en röd boll och en tjej som står framför med en tigerskjorta.
En bicyklist som hoppar med sin cykel i luften
En blond kvinna håller ett föremål i munnen och en rosa tandborste i handen medan hon sitter framför en färgstark soffa.
Två personer på toppen av en klippa
Den svarta hunden är i vattnet på stranden.
En pojke gör en tå beröring framför ett träd.
En man som klättrar uppför ett berg.
En liten pojke springer runt medan andra tittar på en scen.
En gammal kvinna i svart klänning håller en limpa bröd utanför en dörr.
Folk som går runt i centrum av en stad.
Fyra män hänger framför en byggnad.
En kvinna i en rosa blus samtalar med en road manlig kaukasier.
En man i svart väst och färgstark slips drar uppmärksamheten till en publik nära en uteservering.
En ung kvinna vilar huvudet på en mans axel.
En äldre kvinna i flera lager kläder stickar ett plagg som, hon sitter nära en uppsättning trappor.
En man som bär på en kvast och en soptunna tittar på medan en ung pojke skiner på en kvinnas sko.
3 män i t-shirt och shorts sitter på gräs äter mat.
Ett barns ben klämmer genom en hunddörr.
Rödskjortad arbetare klättrar stege för att kika in i en behållare uppfälld på en gaffeltruck.
En tjej med blont hår hoppar från en däcksvinge.
En ung kvinna som dansar för en liten publik.
Barn och mammor sitter i halvmåne på golvet.
En gråhårig kvinna vänder sidorna i en bok för en cirkel av barn sitter i blå stolar.
Barn äter vid ett långt bord med svarta stolar.
En kvinna med flätat hår sitter vid ett bord fullt av mat och gerting.
En snowboardåkare använder en ramp för att slipa en räls.
En gul och brun hund går på toaletten utanför.
En man som bär gul rock står på toppen av ett berg.
En stor gentleman vet inte hur han ska använda sitt paraply.
En man som sitter på en stol mitt i en grupp.
En kvinna på en bakgårdsfest hoppar rep på gräset.
En kvinna som sitter vid ett picknickbord håller ett barn.
Män i röda bågar sjunger i en kör.
En pojke hoppar i en pool.
Ett ungt spädbarn i en vit topp som gråter.
En man i blå skjorta som skriver på en krittavla.
En man med grå handskar håller händerna mot öronen på ett trapphus.
En ung man breakdancing på en kullerstensväg med många människor tittar på honom.
En man som går medan han håller en hatt på en pinne.
En brunett kvinna smakar sin ätliga skapelse från en skål.
En stor brun hund springer med ett grönt föremål i munnen
En säkerhetsofficer ser ut över vatten där det finns ljus.
Ett litet barn är med vått hår står vid poolen insvept i en handduk.
Dessa berg paret tittar på våra vackra.
En gentleman i telefonen vid sitt skrivbord medan ett barn sitter i knät och ritar på ett papper
Tjej i rött, med randiga tights, spela fiol utanför byggnaden.
Många svarta hundar springer i ett gräsområde.
En kvinna som ler när hon jobbar med en maskin.
En ung flicka klättrar på klipporna samtidigt som hon är säkert bunden uppifrån.
En ljusbrun hund petar in huvudet i borsten.
En man och en kvinna går förbi bänkar med utsikt över vattnet.
En tennisspelare som rör sig för att träffa den annalkande tennisbollen.
En man i grå skjorta och svarta byxor spelar tennis.
En ung dam tränar tennis.
Manlig barn spela på runda inneslutna rida i parken själv.
En kvinna på ett café dricker kaffe medan hon gör pappersarbete.
En person i röd hatt som bär på en stor skål med glass med flera kottar som stinker av den.
Tre kvinnor sitter runt en upphöjd eldgruva och kokar stekta smågrisar.
En person håller i en cykel i luften med sin kropp i flygläge.
Två män pratar med varandra medan de sitter vid ett bord, och en håller i en delvis öppen bok.
En man med röd hatt sitter på en pall på sidan av vägen.
En hund sträcker sig över det bruna gräset.
En man gör en backflip medan han försöker hoppa på en cykel.
En bebis i en grön väska kikar ut.
En man med grått hår sätter en svart krage skjorta över en vit knapp-up skjorta medan flera andra män tittar.
Ett band spelar badat i scenljus.
En man i svart jacka spelar en svart elgitarr och sjunger.
En leende person med en färgstark mohawk frisyr.
En stor vit pudel går på gräset och bär en sandal.
Två flickor håller upp sin yngre syster.
En man i en kilt spelar ett instrument framför en butiksfront.
En liten pojke dricker vatten från den gröna slangen.
En kvinna cyklar nerför en trottoar, när män i långa kostymrockar står runt med en rad andra människor.
En ensam surfare som rider en enorm våg i havet.
En pojke med orange skjorta har håret rakt upp från huvudet.
En ung flicka i rosa klänning stirrar på en tunnelbanetidning rack.
Två personer står i grunt vatten och viftar med gnistor
Två kvinnor i ett jordbrukslandskap som sorterar grödor.
En man på en fyrhjuling hoppar på ett fält.
Kvinnor som cyklar moped och motorcykel.
En dam håller ett paraply bakom vad som också ser ut att vara ett vattenfall.
En man och en kvinna som står vid en disk med mat.
En cowboy står nära två får och en hund på en rodeo.
Tre män utomhus ler, dricker öl och tar bilder.
En ung kvinna i en tanktopp röker en cigarett medan hon håller i två boccebollar.
Några personer på en kanot i vattnet.
En man med dreadlocks ler medan han sitter i ett dj-bås.
En man häller något i en kopp från en dryckesmaskin.
En man som bär en skjorta som säger "pengar pratar" är att dricka vatten medan luta sig mot en Verizon lastbil.
En stor brun hund sniffar en liten vit hunds bak.
Två blonda flickor i vita klänningar, den ena mycket mindre än den andra, står på stranden av en stor vattenförekomst.
En man med arm runt flickvännens axel när de tittar på något.
En man sitter inne i en brevlåda med en telefon i handen.
En svart hund är i en hundkapplöpning.
Två kvinnor står bredvid varandra och skrattar.
En flicka och hennes barn går bredvid ett berg.
En man i vit t-shirt och beige shorts sover på en svart soffa.
En ung pojke pekar och tittar på ett träd med fler träd i bakgrunden.
En liten svart pojke i blå skjorta och mörka shorts som springer genom en fontän.
Folk som har kul på en grillfest.
Två vuxna och ett barn står på en klippa med berg i bakgrunden.
En ung man i t-shirt ler i en bokhandel.
En grupp män som bär hjälm står i en linje med flaggor och en publik i bakgrunden.
En orange lastbil kör nerför gatan framför en vit byggnad.
En baseballspelare står på plats och fångar en flygande baseball i sin handske.
Mannen arbetar efter mörkrets inbrott på en marknad.
En hund vilar på en madrass medan en gammal kvinna sitter på golvet.
En ung pojke leker med en slinky på gatan
En person seglar i luften med en röd fallskärm över gräs.
Män i traditionella skotska kläder marscherar och spelar säckpipa.
En grupp soldater marscherar i led medan de håller flaggor.
Fyra pojkar springer iväg med en lutning.
Två lag av pojkar som spelar fotboll och en pojke är uppe i luften med bollen bakom sig.
Ett barn som leker med vattennudlar i en pool.
En tjej i en svart utstyrsel hula hoops medan folk sitter vid borden och äter.
En person står på en klippa med utsikt över en bred dalgång.
Två unga pojkar sitter i en stol med blommor och en grön kratta.
En fem mans övningsteam på scenen.
En brud och brudgummen småpratar med en gäst när brudgummen skakar gästens hand.
Par som är gifta i en kyrka.
Två personer rider ner en stock flume i en nöjespark.
Två unga män deltar i en fotbollsmatch.
Den här killen är i luften när han bär en röd fotbollsuniform.
En kvinna som lagar mat på spisen.
En tjej med svarta handskar springer.
En tjej i blå jeans lutar sig mot en guldgul bil.
En man och en pojke poserar för en bild i en trappa med utsikt över ett vattenfall.
En kvinna med lila jacka står bredvid en häst.
En brud kramar en person med kort blont hår.
En rödhårig kvinna med gröna ögon går in i en skåpbil.
En man i en rutig skjorta står nära en hög med spillror.
Barn leker med en cykel i sanden.
Tre små pojkar brottas och en är skjortlös, leende, och vänd mot kameran.
Pojke i orange, hoppa från en rostig färgad pipa, i sand.
Två män i grå skjortor och röda hattar arbetar med cement.
En kille som tar en tupplur i baksätet på ett fordon.
Fordon parkerade på en restaurang och bensinstation någonstans i Mexiko.
Två flickor är i kö för att beställa på ett mexikanskt matställe.
En vän foto med två pojkar tittar på varandra medan flickan tittar på kameran leende.
En svart och brun hund vilar huvudet på nedre trappan.
En liten pojke i röd skjorta som svingar ett basebollträ
Man i affärskläder hoppar från sidan av en byggnad.
Två män sover i baksätet på en bil.
Ett par i bilen tittar på något bortom kameran.
En kvinna klädd i svart och rosa har en stor tatuering på ryggen.
Två killar som ler när de sitter i ett fordon.
Män och kvinnor cyklar i en varm solig dag i en stor stad.
En pojke i gul tanktopp som skrattar på en strand.
Ett par sitter på en skuggad bänk med utsikt över träd och en stor byggnad.
En infödd pojke, i gult, svänger från ett rep.
En grupp barn leker i vatten.
En grupp människor springer på sanden.
Walkers och cyklists beger sig ner på en tom New York-gata.
Man håller en liten flicka på en gata.
En våt ung flicka i vit rock står bland vattenfontäner.
Två honor blåser bubblor med sitt tuggummi.
En vuxen man och ett litet barn tittar till vänster när de cyklar.
En vit bil står parkerad bredvid några hus i ett tredje land.
Fem män bygger en grund för ett hus
Ett barn simmar under vattnet i en pool.
En man som bär röd hatt medan han håller i en stege med en man i brun hatt och tittar på honom.
Två barn jagar varandra i sanden.
En grupp människor som tittar över räcket på vattnet och marken täckt av dimma.
En grupp människor plockar grönsaker utanför.
En man lyssnar på någon i telefonen med en främmande blick i ansiktet bakom ett fruktstånd.
Vuxna och barn som går på en grusväg.
En person i blått undersöker en vägg.
Män arbetar tillsammans med ett byggprojekt.
En person med randiga röda strumpor springer på en skogsväg på kullen.
Folk på gatan går förbi en dockteater.
En brun hund som bär munkorg springer på sand.
En pojke med röd skjorta och blå shorts går ut.
En man i blå skjorta och grå byxor sover på en trottoarbänk.
Byggarbetare bygger en ram för en struktur.
En grupp människor bygger en mur för en byggnad.
En kvinna spelar orgeln i en kyrka.
En ung man i en keps spelar elgitarr.
Män som arbetar med konstruktion håller upp ramen för en vägg.
En man i svart rock äter en munk medan andra män ser ur bild.
Fyra personer står framför träd.
En man med mohawk frisyr bär en ryggsäck på ett college campus.
Två barn glider i snön.
En brindle hund springer bredvid några pålar i marken vid vattensidan.
En man är utanför och säljer olika leksaker.
Kvinnan i den gröna randiga skjortan och ryggsäcken har en tatuering på ryggen.
En gatuartist rider en hög enhjuling samtidigt balansera jonglering enheter.
Fyra män och en kvinna som sitter på marken i skuggan.
Hunden springer genom djup snö.
En man jobbar på kaboosen på det röda tåget.
Den lille pojken springer genom sprinklern.
En grupp människor bygger en ram av en byggnad.
En person tittar på vattenstrålar.
En man ligger på två gröna luftmadrasser med en tumme upp.
En man med huva som arbetar i en kiosk visar upp sina varor.
En vy över en marknadsplats full av människor i ett asiskt land.
En man som står i sitt nät fiskar i vattnet.
Två män i vita t-shirts och verktygsbälten sitter på ramarbete för en struktur.
En grupp människor äter en måltid utomhus tillsammans.
Tre personer får sin bild tagen när en är böjd över.
De tre hundarna står i sanden.
En flicka är på väg ut ur en simbassäng.
Människor som ligger och sitter nära viss ljud- och visuell utrustning.
Flera personer är i en byggnad med luftmadrasser och andra tillhörigheter.
Pojken och flickan bär simglasögon.
Här är en bild på ett barn klädd i kostym, leende och dans.
En mor, klädd i traditionella kläder, och hennes två barn poserar för en bild.
En motorcykelförare kör en svart motorcykel.
Flera unga pojkar och flickor hoppar på en studsmatta utomhus.
En dam med mörkt hår som tittar på några papper på tunnelbanestationen.
Två vandrare står på toppen av ett snöigt berg.
Man och kvinnor som tittar på ett paket en frukt på en livsmedelsmarknad.
En svart hund hoppar över en stolpe på grönt gräs.
En dam som sitter bredvid en Sprite-flaska och slickar något vitt på gaffeln.
Den skadade idrottsmannen bärs av flera personer.
Ett litet barn hoppar upp i luften ovanför havet.
En hund simmar i vattnet.
En skara människor på en mässa ser tre män reta upp en stor tjur.
En läkare på ett kontor som ler mot kameran.
En man och en gammal kvinna står och tittar på något bakom fotografen.
Ett paraply som skuggar en ung kvinna med en liten pojke som hukar sig under bordet.
En flicka är på väg att sparka en fotboll i gräset.
En tjur som anfaller en tjurryttare i en live rodeo.
En svart man i en svart dräkt står framför ett tunnelbanetåg.
En pojke som spelar på ett arrangemang av stenar.
En liten pojke som bär en ljusblå skjorta ler när han håller något i handen.
En kvinna i baddräkt går en hund på stranden.
En kvinna i en butik med gula ballonger.
Kvinnan läser en bok.
Två flickor som ligger i gräset ler när deras bild är tagen.
Killen med skidjacka hoppar från bron i vattnet
Fem män står utanför och ser ut som om de är på väg att arbeta.
En man i orange jacka pratar med en kassörska.
En blond tjej i rosa baddräkt som springer genom sprinklern.
De två unga pojken äter mat.
Tre vuxna och tre barn simmar i en allmän pool med ett barn redo att dyka.
En person på en cykel rider genom ett skogsområde.
Ett barn i orange är på en boogietavla i vågorna.
En dam i blått, tar en närmare titt på omgivningen genom att titta i stående kameran på parken.
Bilder på en vit tegelvägg med en leende man som står framför väggen.
Folk går på kakel på en utomhusmarknad.
En man i grön skjorta och svarta byxor tittar in i en affär på en fullsatt marknadsgata.
Ett gäng shoppare som tittar på TV-skärmarna i en butik.
En greyhoundhund springer runt ett spår.
Tre barn på dykbräda, med ett hoppande av.
Två äldre kvinnor sitter på en vit bänk i en park.
En grupp människor väntar i kön för ett spel.
Tre män klädda som kockar sitter på en stenbänk.
En man som går ut ur ett portabelt badrum.
En liten pojke i vit skjorta och jeans stoppar fingrarna i munnen.
En hund som springer genom sanden.
En man och en kvinna omfamnar medan de står mot ett grönt Heineken-tecken.
Brunhårig man med en vit skjorta som visar upp ett leende med öppna armar.
Ett barn ligger på en handduk och gråter när de byter blöja.
Två män som ler framför en eldsvåda.
Flera asiatiska kvinnor klädda i svarta kläder och kronor håller tallrikar med mat på dem.
Folk hoppar fallskärm.
En person ligger i vattnet och kastar tillbaka håret.
Ung skäggig man som bär en vit tanktopp sitter bakom ett trumset.
En svart hund hoppar i luften medan en kvinna skriker i bakgrunden.
Många barn i elementär ålder samlades och satt utomhus.
Två pojkar i shorts sitter med en surfplatta med andra människor i bakgrunden.
En svart och vit hund springer genom gräset.
En man som spelar gitarr i ett sovrum med en svampbild på väggen bakom sig.
En blond kvinna lämnar en röd stolpe.
En liten pojke i grön overall kastar upp händerna bakom det blanka restaurangbordet.
En välklädd flintskallig man med röda glasögon går i full fart.
Olika människor köper, och tittar på olika typer av grönsaker och blommor.
En flicka i gul skjorta sprutar två personer med vatten.
En liten flicka hoppar ner från dykbordet i en pool.
Tjejen skriker med rosetter i håret.
Ung man visar sin tunga piercing medan en kvinna står bredvid honom
En simmare simmar över en knäpool.
En man i blå skjorta som ger sitt barn en klunk av sin drink.
En kvinna i ett rum justerar hängande kläder.
En gentleman med bruna byxor och skjorta pratar med en man med vit skjorta framför en symaskin.
En utklädd kvinna spelar ett instrument på en bänk.
En kvinna, i en röd baddräkt, justerar sina simglasögon medan hon står vid en pool.
Två små barn leker med leksaker.
En kvinna använder en tidning för att ge skugga och bli av med bländning medan hon använder sin dator utanför.
En skateboardåkare utför ett skateboardtrick mot en graffitivägg.
En ung pojke, som bär en röd fotbollströja, strumpor och klapperskor, står på ett fält av grönt gräs.
Mannen sitter på en grön stol med fiskespö i vattnet
En blond pojke i en mörk huva håller i ett fiskespö.
Två personer forsar nerför en flod nära tallar.
Två personer paddlar en kanot nerför en grov flodsträcka nära en tallskog.
En pojke hoppar ner i vattnet påklädd.
En turistbuss fullpackad med människor när de alla tittar åt vänster, anstränger ögonen på ett ämne som guiden påpekade.
En kvinna håller i en annan kvinnas arm.
En vit hund bär en boll över gräset i närheten ett staket.
En man i gul jacka åker skidor i snön.
En saxofonspelare klädd i en blå tröja och en dragspelsspelare underhåller människor på gatan, inklusive en pirat.
En indisk man som står på stranden av en flod.
Gult lag mot rött lag sparkar en blå &amp; vit fotboll.
En liten pojke närmar sig fotbollen för att sparka den.
En man med skägg och solglasögon lutar sig tillbaka på en soffa med fötterna på ett soffbord.
Ett barn i rosa kläder stirrar på majs på kokset
Ett barn som är täckt av en vit filt sover.
En pappa firar en födelsedag med sin familj via webcam.
Tre män och en kvinna hoppar in i en pool full av lugnt blått vatten.
En brun hund som jagas på landsbygden
En gift brud och brudgum som går längs trottoaren och har ett intimt ögonblick.
Dam klädd i en exotisk klänning.
En kille i strippskjorta som ligger på en picknickfilt och tar en tupplur.
Två män förbereder jorden för plantering av nya grödor.
En gråhårig kvinna i gul skjorta som sitter under ett blått tecken.
Det finns en stor grupp människor på scenen som håller flaggor.
Den här pojken sprider armarna medan han leker i vattnet.
Ett ungt par som stirrar framför havet.
En ung kvinna med långt brunt hår, spelar en svart gitarr, vänsterhänt.
En weiner hund fångar en blå och gul tennisboll.
En man går på gatan med solglasögon på huvudet.
Två personer står mot en vägg efter ett träningspass.
En häst hoppar två räcken med en ryttare i grön jacka.
En man står bredvid en svart fällbar stol.
Fem personer vadar och simmar vid kanten av en flod eller sjö.
En man använder sin säljtelefon nära några hängande mattor.
Det sitter en tonårspojke i något som verkar vara någon sortsrickshaw, medan föraren pekar på honom bakifrån.
En flintskallig man sitter på trottoaren lutad mot ett gäng vävda filtar.
En ung kvinna i svart bikini borstar sitt långa bruna hår på stranden.
Ungt barn plaskar och leker på stranden.
En man i vit skjorta och grå byxor arbetar i en klädaffär utomhus.
Sidewalk försäljare klädd i vit skjorta bruna byxor säljer grillad majs.
En hane och två honor (båda i baddräkter) står bredvid ett sandslott på stranden.
En man som ser ut som en staty på trottoaren.
En man i en grå tanktopp med halmhatt som sjunger till en mikrofon som spelar gitarr.
En man står framför ett bildspel och ger en presentation.
En ung flicka i en rosa bikini skrattar längst ner i en vattenrutschbana.
Den bruna hunden springer genom ett fält, med en boll i munnen.
En ung pojke i vit skjorta med gummiklubba.
Flicka i klänning hängande på orange räcken
En grupp vuxna som håller i musikinstrument verkar inte spela på instrumenten.
Folk som sitter ute på grönt gräs.
Barn skriker och går över sand, en annan figur och havet i bakgrunden.
Man sprutar volleyboll över nätet med en annan spelare framför sig.
4 stränginstrument som spelar män sitter på en svart scen och spelar sina instrument från deras musikställningar.
En man i en stockrock som kantar marken.
Två österländska män klädda i vita dräkter spelar en stor gitarr och en bongo.
En riddare på hästryggen och en annan man återuppväcker en medeltida scen för en grupp åskådare.
Två unga flickor hoppar av eller över en betongbarriär i en innerstadspark.
En kvinna i randig tröja står på en kulle.
En äldre man i blå kostym går ut ur en byggnad med namnet "Grace" på framsidan av den.
Den svarta hunden hoppar upp ur vattnet med något i munnen.
En leende pojke hänger på en zip-line struktur på en lekplats.
En grupp poliser utanför en stadsbyggnad.
En man i en blå kula och utan skjorta som arbetar på ett tak.
En grupp människor omgivna av träd, ta en hötur tillsammans i solskenet.
En man med glasögon kysser en kvinna i pannan.
En vigselceremoni i en kyrka.
En kvinna med axellångt hår sitter på en trottoar med en blå randig skjorta och höga klackar.
En blondhårig kvinna sitter bredvid en hög ryggsäckar.
En grupp orientaliska dansare uppträder på en parkeringsplats.
Två små bruna och vita hundar står tillsammans.
En man och en kvinna ligger på knä framför gången och gifter sig.
En ringbärare som bär en ringklocka på en kudde på ett bröllop.
Tre unga män spelar ett spel av Monopol där två av dem fysiskt argumenterar.
En hund som sniffar på borstarna medan en tjur tittar på
Två män och en kvinna står tillsammans på en våt gata med jackor, hattar, och kvinnan bär ett paraply.
En kvinna viftar med handen från ett fönster.
En kvinna i brun skjorta och en tiara pratar i telefon.
En polis i en skinnjacka står vid sin motorcykel.
En vit hund springer mot kameran.
En man på en gräsklippare kör förbi en bil.
Blond man med vit knapp upp skjorta framför två rödhåriga kvinnor, en använder en mikrofon den andra bär hörlurar.
Den här personen bär en svetsmask.
En överviktig man bär en skyddande hatt och handskar.
En vuxen som spelar schack med en ung blondhårig pojke.
Tre svarta hundar är på en strand.
En läkare kontrollerar en ung flickas hjärtslag.
En grupp barn står i rad och håller pinnar och svärd.
En kvinna piskar upp håret ur vattnet.
Ett band av fyra gitarrister och en trummis uppträder på scenen.
Det är en konsert på gång.
En casinoåterförsäljare och ett par ler mot kameran.
En man med blå hjälm är på en motorcykel.
En rödhårig clown gråter tårar i en vit hatt på scenen.
En kvinna i vitt gör akrobatik.
Två personer är klädda i "leotards" som uppträder.
En ung pojke som hoppar från en lekplatsleksak.
Den lille pojken som bär den blå skjortan äter med ätpinnar.
En Budweiser-sponsrad racerbil accelererar snabbt med rök bakom sig.
Man på en lång enhjuling, som bär ljusgul skjorta, röd bandanna och kamouflage byxor jonglerar 3 stift medan folk tittar.
En gammal kvinna i en halsduk är i stan.
Ett barn bär en pappershatt och äter på ett matställe.
En svart och vit hund hoppar för en tennisboll.
Två hundar som bär tävlingsutrustning springer på lerig mark.
Tre killar är mitt uppe i backflips.
En spelare sparkar fotbollen från hörnet av fältet.
Bmx MC Hoppar av rampen
En pojke försöker hålla balansen medan han står på två flytande apparater medan två andra tittar.
Man pekar på en kvinna som sitter ner för att äta.
Två män står framför kassaapparaten med flera saker.
En kvinna i vit skjorta bär glasögon.
En fönstertvätt i en blå skjorta tvålar upp fönstren.
Två människor här bär något runt halsen.
En grupp kvinnor i vita dräkter går genom gräset.
Person som håller en gitarr med religiösa bilder och reflekterande klistermärken på framsidan.
Två män står framför en protestskylt på en röd elektrisk låda.
Flera män och kvinnor njuter av mat utomhus.
En kvinna med randig topp står nära uppstoppade djurpriser.
En blond tjej spelar på en uppblåst hoppleksak.
En man i vit t-shirt tittar på en hund gör en backflip
Killen i randig skjorta spelar sin elgitarr.
En kvinna tränar gymnastik medan en man fotograferar henne i luften.
En stolpevalvare är på väg att avfyras från golvet med sin stolpe.
En man i halmhatt gräver med en spade.
En kvinna med rött hår håller i två katter.
En pojke klädd i grönt rider en video motorcykel spel framför skidboll maskiner.
Två kvinnor spelar volleyboll på sanden.
Damen har en vacker vit klänning ihopkopplad med en vacker vit högklackade skor.
En liten pojke som står i mycket högt grönt gräs.
En man hanterar sin nästan tomma drink medan han skrattar åt något på andra sidan bordet.
En fotbollsspelare springer på planen
En flicka i röd skjorta färger som hon står vid sitt skrivbord.
En ung pojke öppnar en present.
Ett barn med blå skjorta och blå byxor står i en park.
En ung pojke som står mellan en vägg och flera stora stenblock.
En flock hundar springer iväg längs ett spår.
En flygkvinna kollar en äldre kvinna.
En grupp män klädda som pirater står utanför Cheesecake Factory med skyltar.
En ung pojke skriker på en berg-och dalbana.
En man klädd som en indian med två hundar som står och pratar med en grupp människor med lite hö.
En kvinna skriver en lapp för en äldre kvinna.
En vältränad volleybollspelare förbereder sig för en gupp.
En man tittar ut genom träbarer, som han håller i sina händer.
Närbild av bartender (kvinnor) ta tag i ett glas i baren.
Man och pojke med ryggsäckar på en vandringsled.
En hund springer på en gård med en deflaterad boll i munnen.
Flickan återfår lugnet i en solnedgång med en man i bakgrunden
På natten sitter en ung man nära ett bord som innehåller aluminiumfolie, choklad och kex.
Två män steker marshmallows utanför vid en lägereld.
En kvinna i en ko mönstrad förkläde och faux ost topp hatt skär riktig ost.
En brun och vit hund tittar in i en pool på en tennisboll.
En man i orange skyddsväst vänder sig till flera andra män i en skog.
En hejarklackstrupp poserar för en bild framför fullt blekmedel
En liten vit hund har koppel och går bredvid ett staket.
En man använder en motorsåg för att rista en träskulptur.
Tre nyhetsutgivare, två män och en kvinna, sitter vid nyhetsdisken och skrattar.
Pojken i röda glasögon simmar under vattnet.
En liten, leende pojke i en blå skyddshjälm och gul skjorta rider sin skoter på en trottoar.
Två hundar antingen slåss eller leker tillsammans.
Ett litet barn som bär blå topp är på en blå leksak.
En grupp människor i baddräkt poserar för en bild.
En liten pojke med brunt hår hoppade ner från en brun stol på golvet.
Pojken bär badbyxor håller goggles och löpning
Barn som leker med en hulahoop på en cementuppfart i bostäder mycket.
Folk går upp för en rulltrappa i köpcentret.
En liten pojke i grön skjorta begravs upp till midjan i sand.
En kvinna i orange jacka pratar på sin mobil.
En kvinna serverar en kopp soppa från en stor gryta med soppa.
En man med hatt bygger ett hus.
Någon i en blå skjorta som skriver på en del av en tidning.
En hund försöker dricka vatten från en sprinkler.
Män i hårda hattar som arbetar med en stor guldmaskin som utför vägarbete.
En gammal man cyklar på en landsväg.
En pojke i en gul tank topp springer bort från en kraschande våg.
En man i blå skjorta som tar en bild av ett berg.
Här är en bild av elever i ett klassrum som gör ett datortest.
Ett barn som bär hatt står på en strand och tittar ut över havet.
Ett litet barn klättrar upp för en röd matta på en festlig matta.
Man med orange hård hatt, kör ett byggnadsfordon och vinkar.
En man som bär en bygghatt och väst går framför en stoppad stor röd semi i ett skogsområde.
Man skjuter bilder på kvinnor på stranden.
En man som bär glasögon och en grön skjorta övar spela ett stränginstrument inomhus.
Två små pojkar som cyklar på gatan.
Barn med shorts som leker utomhus i parken med sprinklervatten.
En brun hund bär en våt pinne på havets strand.
Två män i fåniga glasögon sitter på golvet.
Två byggnadsarbetare sitter på några rör medan en vågor, dunkel hans ansikte.
Människor som sitter vid långa bord alla vända åt samma håll, en del skrivande och en del tittande.
En man och en kvinna som hoppar från en båt i blått vatten.
En kvinnlig softballspelare glider dramatiskt in i en platta när basmannen står redo att fånga bollen.
En flicka öppnar en present medan en ung pojke i blå pyjamas klockor.
Två hundar hoppar upp mot varandra på ett gräsfält.
En pojke går genom en parkeringsplats fylld med bilar.
En man i brun läderväst och en kvinna klädd i rött och svart som håller om varandra.
Folk i en auditorium väntar på att något ska börja.
En person som bär jeans sitter ovanpå en hästsadel.
En underhållsarbetare klättrar in i sin gröna lastbil.
En man med svart hår och brun skjorta skapar porträtt av människor.
Mannen bär glasögon och en grön skjorta, utför en uppgift på en dator.
En närbild av en liten pojke som ler samtidigt som han håller fast vid någon lekplatsutrustning.
En kvinna bär på en ung pojke medan hon skrattar med en man i grå t-shirt.
En mormor tittar på sin dotter och sonson leka med tåg i ett vardagsrum.
En ung hane dricker på en juice.
En kvinnlig sångare sjunger passionerat medan back-up gitarristen spelar i bakgrunden.
Människor står på toppen av en röd turistbuss
Ett litet barn springer längs en strand när fåglar flyger bland honom.
En liten hund fångar en tennisboll i munnen.
En polis står utanför på gatan med händerna i fickorna.
En person i ett fält tittar genom ett teleskop medan en blå bil närmar sig eller väntar.
Fordonet korsar en vattenström i ett skogsområde.
En man som bär Jean flyger en drake nära stranden.
En ung man som slappnar av sina ben på en pice av maskiner
Två unga flickor ler och skrattar.
En man i rosa t-shirt sjunger en sång
Någon matar en jordgubb med en sköldpadda.
Hunden hoppar över de höga hoppstängerna i en hundshow som ägaren tittar på.
En hund på en tävling kör ner en ramp.
Hunden springer runt en vit och rosa stolpe.
En vit kärra som kör en racerbana.
En grupp barn leker i vattenfontänen.
Sex små flickor sitter på en cement kulle.
En liten pojke i en mörk t-shirt och jeans tar stor glädje stående nära en fontän utomhus.
En långhårig kille som gör en backflip på studsmattan.
En person i en randig fleece klipper en karbiner på en metalllinje.
En bil är i vattnet
En man sitter på en hög mattor vid en byggnad medan ytterligare tre män och en kvinna står i närheten.
En man skateboardar och en annan nan hoppar över hans huvud.
Fyra unga flickor som leker i vattnet.
Två män och en kvinna sitter på en bänk med en clown.
En pojke och en man som verkar vara pojkarnas far arbetar med ett konstprojekt tillsammans.
En äldre man gör sig redo att klippa sig hos en frisör.
En äldre man sitter vid en arbetsbänk medan han ristar sin konst.
En ung munk i rött och orange sveper golvet.
En kille med röd rock, vita jodhpurs och svarta stövlar hoppar sin grå häst över stolpar under en brant tävling.
En vandrare klättrar uppför en stenig kulle med dimma omger honom.
En ung man i glas dricker öl och håller klöver tio i pannan.
Två barn tittar ner och klämmer genom ett stängsel.
Den korthåriga hunden springer över en gräsbevuxen gård.
En hund som springer längs en grusväg.
En liten flicka sitter vid ett bord utomhus och äter vattenmelon.
Tre kvinnor på gatan med träd i bakgrunden.
En grupp människor står i smutsen nära två stationsvagnar, med några säckar på baksidan av en stationsvagn och andra säckar staplade på jorden.
Människor står på en strand, en under ett grönt paraply
Den svarta hunden fångar en leksak i munnen medan han springer ut på fältet.
Två personer väntar på en busshållplats.
Det finns en kvinna, flera män och flera barn på en trottoar där man säljer produkter.
En ung man sitter på en soffa och röker.
En ung man som bär hatt och träningsoverall sitter i förarsätet i en liten taxi.
Tre personer, bogserade av dem kvinnor, är på en strand klädda i tillfälliga sommarkläder.
En kvinna lagar mat i affären.
En ung kvinna håller sin väns cykel åt honom medan han drar ut sin skateboard.
En arbetare korsar bjälkarna i en byggnad som håller på att byggas.
Två män talar i en klubb med gröna gardiner.
En ung man och kvinna både i bruna skjortor sitter och skrattar.
En kvinna i röd klänning som spelar ett instrument.
En kvinna sitter på stranden täckt av mycket sjögräs.
En pojke på sin cykel stannar och tittar tillbaka på kameramannen.
Detta är en kvinna i gul rock som letar efter något hon tappade medan hennes manliga följeslagare stirrar på kameran.
Två barn rider på en nöjespark.
Två olyckliga äldre människor som tittar förbi kameran, mannen som håller i en bok och kvinnan som bär päls.
En man sitter med foten på en stolpe och ler.
En svart och vit hund bär en vit frisbee över gräset.
Skolförsäljning för att tjäna pengar på resor.
Ung flicka bär rosa hatt och jacka och blå skjorta hoppa i pölar
Mannen tränar en hund att sicksacka genom stolpar.
En skallig man i röd skjorta uppträder framför en folkmassa.
En kvinna med tatuering spelar saxofon.
Folk sitter och kopplar av bredvid en pool i en plaza.
Person i silhuett tar en bild av en stor klocka.
Två kvinnor köper en produkt som den ena kvinnan i den gröna toboggan säljer.
En ung pojke i blå skjorta leker med en leksaksbil.
Tre vita barn leker med LEGO och leksaksbilar på mattan.
Mamman ser sitt barn leka med solglasögonen vid fönstret.
Två små pojkar delar en baby sving i skymningen.
En kaukasisk man och hans son som hade tid att umgås.
En fotbollsspelare, hans hjälm halvvägs, tittar på marken.
Den lille pojken är på väg att gå in i sprinklern.
Två hundar, en brun och den andra svart, leker i surfingen i det grunda havsvattnet.
En man ses hosta på en fullsatt gata.
En brun hund hoppar över en lila och grön grind.
En fotbollsspelare förbereder sig för att kasta bollen.
Folk ser på när en hund skalar en trävägg på ett gräsfält.
En Elton John ser ut som en kille som spelar ett instrument på scenen.
En man och en kvinna som dansar framför målningar hängande på en vägg.
Ett barn förbereder sig för att kämpa med en karneval attraktion.
I en stor stad samlades många människor runt ett stort reflekterande ovalt konstverk.
Graffiti täcker de flesta öppna ytorna i den här bilden.
En man utan skjorta klättrar på en klippavsats.
En stor grupp människor är på en strand.
En man som går längs en väg bredvid en blå byggnad och röd stoppskylt.
En hund leker fånga på grässlätten
En kvinna öppnar en gåva medan hon står i en matsal som är festligt dekorerad: hennes ansikte hindras av en av dekorationerna.
En liten hund leker med en färgglad boll i sanden.
En svart och vit hund som hoppar i luften för att fånga en vit frisbee.
Svart hund hoppar upp i luften för att fånga en frisbee.
Två barn i kampsportskläder slåss på en blå matta.
En tjej som klättrar upp i ett rockansikte.
Gammal kvinna i vit hatt sitter på en låda och tittar på skjortor på ett bord.
Arbetare reparerar en del av vägen.
En man med grå mössa, guldsmycken och vinterkläder tittar på något i fjärran.
En orange båt lämnar stranden medan en person tittar i närheten.
En man med svart mustasch skär kött med en stor kniv.
En man på toppen av en häst som ler mot kameran nedanför ett berg.
En pojke i blå skjorta och glasögon står vid ett träd.
Underhållningsgäster vid en renässansfest som bevakas av åskådare.
En man skriker åt någon från ett spelbås.
En man med solglasögon i rosa skjorta.
En kvinna skriver i en dagbok, medan hon sitter på en bänk på ett kafé.
Två pudlar som leker med en röd leksak.
Två män inspekterar och fixerar däcket på en röd inramad, gul kluven cykel med cykelstolen mot marken.
En person surfar på en våg medan en annan person går mot den.
En ung man som bär AIDS WALK t-shirt står och skriver på laptopen.
En man klädd i svart står med tre kvinnor som har blont hår.
Två bruna hundar leker i ett snöigt fält.
Ett barn leker i en pool medan det bär orange floaties.
En ung pojke och en äldre kvinna som sitter vid ett brunt bord i ett blått rum.
En man och kvinnor är ute på Farmosa och tittar på menyer när de chattar.
Det finns en man som bär röd skjorta och bruna shorts hoppar upp för att slå en tennisboll med en racket.
Fyra småbarn underhålls av en dragspelsspelare.
Två kvinnor som sitter under ett L.E.D. tecken på en person som går.
En man som står utanför en affär på gatan.
Två personer står armbåge djupt i havet och tittar på solnedgången.
Tre pojkar leker i en ofullbordad byggnad.
En ung pojke verkar hamra metall ovanpå ett städ.
En kvinna, som bär halmhatt, presenterar en mängd olika varor.
Den vita och bruna hunden springer genom gräset.
En tjej i röd jacka skrattar åt kameran.
En kvinna i blommig klänning går nerför gatan förbi sin spegelbild.
En man i randig skjorta som hackar svamp.
En person som klättrar på en sten medan andra står och tittar på.
Männen i Gators hjälmar har sina armar lindade runt varandra.
En skjortlös man jobbar på ett tak.
En grupp människor på en olympisk händelse.
En man i en gul regnrock viftar med den kinesiska flaggan under en regnig händelse.
Folk som står på sand i regnet.
En asiatisk idrottsman i en ljus jacka ifrågasätts av många reportrar som bär regnjackor.
En folkskara samlas runt en kvinna som spänner sitt huvud
Tre personer står framför en skylt från Peking 2008.
En man med hatt tar ett foto med kameran, medan en förbipasserande ser irriterad ut.
En grupp människor står i ett rum med takfönster.
En blond kvinna har ett paraply över en racerförare.
Två äldre män arbetar för att reparera ett stenstaket nära en stuga.
En man bär hatt och vit skjorta.
Ett gift par går upp för trapporna.
Man med t-shirt och khaki shorts knäböjer på marken.
En man serverar en volleyboll på sandbanan i en volleybolltävling.
En grupp människor håller upp tre fingrar.
En kvinna som står i en röd bikini på en utomhus sandvolleybollbana.
Flickor i röda bikinin gör en dansrutin på OS 2008.
Människor i kostym och hattar poserar med amerikanska flaggor och fingrar som hålls upp med nummer tre.
Ett barn i röd skjorta klättrar på lekredskap.
En mörkhyad ung flicka får sina gympaskor polerade av en skoputsande pojke i Indien.
Brandbilslinje på båda sidor om en trafikerad tvåvägsväg.
En person som bär Rollerblades hoppar över en gul grind.
En brun hund som gräver efter en boll i sanden
Bild på en röd vagn och en liten pojke som cyklar framför en tegelbyggnad.
Kvinnan håller sin son på de livliga gatorna.
En dam och två små barn sitter på en parkbänk med duvor vid sina fötter.
Vuxna och barn flolic på stranden av en strand.
En grupp människor som bär något inlindat i en amerikansk flagga.
En hund ligger på en madrass på verandan.
Ett par, en man och en kvinna, sitter på en klippa och tittar på havet.
Barn med simglasögon med ansiktet nedsänkt halvvägs
En man i vit kostym går nerför gatan och håller i en tidning.
En lantbrukare gödslar sin trädgård med gödsel med häst och vagn.
Den svarta och bruna hunden hoppar upp i luften för att fånga bollen.
Barn som spelar med en fotboll nära ett målnät.
Flickan simmar med bara huvudet ovanför vattnet.
Två män på hästar jagar ett djur på en rodeo.
Fem kvinnor i klänningar som står i en lobby och pratar.
En man bär en executive klädsel medan han ser något.
Sex män i blå overaller och en man i orange overall går förbi ett varv.
Ungar hoppar på en blå trampolin.
En man paddlar genom några vita vatten.
En kvinna med en kamera ser ut över böljande kullar.
En liten flicka sitter i gräset och balanserar en sten på armen.
En man i röd jacka med jeans på balans i en bowlinghall.
En man med en hink med röd färg märker fisksektioner med siffror.
En man med en penna och papper kontrollera lager.
Två män tittar på kött som står på ett bord medan de antecknar.
Kvinna, med två barn som leker i fontänen utomhus.
En man med keps och shorts sitter på en metallbänk och läser en tidning.
En man i svart skjorta och röd slips som håller i en drink.
En ung man i en blå skjorta som håller en apparat mot munnen och gör en festlig gest.
En vit och svart hund hoppar i vatten.
En man i brun jacka och beigemössa dricker ur en styrofoamkopp.
En kille i svart skjorta hoppar upp i luften på en gångbro.
En man i blå skjorta som hoppar nerför en kulle i en park.
Hund hoppar över röd och vit stolpe medan pojken tittar på
En man som bär solglasögon står framför bandutrustning som håller en gitarr.
En person ligger på gräset med en kundvagn i närheten.
En kvinna som står framför en affär med armarna korsade.
En man och kvinnor som tittar på tidningar i ett fönster.
En pojke i en kedjad gunga ser åt höger och ler.
Ett litet barn sitter medan han håller majs i händerna.
Mannen på cykeln har precis kört igenom lite lera.
Fyra svarta hundar som springer över gräset.
En brun och vit hund går i vatten när man ser tillbaka.
En man kör motorcykel med sin hund i sidvagnen.
Spelare i ett fotbollslag bråkar i ett försök att få bollen.
En liten pojke med blå snopphatt.
Nio män spelar ett spel i parken, skjortor kontra skinn.
Kvinna på salong med svart hår under torkhjälm.
En ung pojke med bara gröna shorts poserar obekvämt med en tegelbakgrund.
Fotbollsspelaren i rött försöker blockera spelaren i vitt.
En ung man i solbränna shorts och grön skjorta faller av sin cykel.
Folk promenerar och samtalar på en trottoar framför ett sjukhus.
En kvinna med en väska pratar med en man på en cykel nära en gata.
En man sitter och gnuggar hakan.
Det finns två ungdomar med ryggsäckar på och sedan står bredvid en vandringsled.
En ung flicka svingar högt med en solnedgång bakom sig.
Två män är i en blå och vit fart båt.
En man och en kvinna i hattar nära en trappa.
Två män med hatt står på den trädklädda trottoaren nära en byggnad.
En hund lägger sig på en stor pinne.
En liten brun och vit hund som fångar en frisbee på en tävling.
En man och hans boskap som kör en vagn på gatan.
En kvinna i sjal håller sitt barn inlindat i en färgglad filt.
En mor och hennes barn poserar för ett foto.
En man kör en grön motorcykel på en våt kapplöpningsbana.
En kvinna håller ett barn och ler.
En man klädd i röd rock, vita byxor och svarta stövlar sitter på en häst på en nöjespark.
En vit rashund som bär nummer åtta löper på banan.
Två män med trasor över ansiktet springer nerför en gata med något som brinner.
Mor och barn på en promenad i en park.
En man på en cykel hoppar över taggiga klippor bland höga tallar.
Två musiker övar för en föreställning.
En överviktig hane spelar elgitarr medan han bär vit hatt.
Kvinnor dyker ner i en swimmingpool.
En flicka tar en bild av sin vän som lutar sig mot ett picknickbord.
En man i hatt jobbar på ett tak.
En man lagar fisk i ett marinblått förkläde.
Två män ser en tredje man grilla kött.
Detta är en natt utsikt över en stad gata med människor och trafik.
Den svarta hunden på fältet har något i munnen.
Mannen med blå skjorta har dreadlocks och solglasögon.
En man i röd skjorta arbetar på en vit skulptur.
De vuxna ler när ett barn leker med några stenar på marken.
En man i orange shorts rör sig riktigt snabbt
En vit hund med röd krage hoppar upp efter en röd frisbee.
Arbetare sågade en stor fisk med en bandsåg.
En man med kort svart hår i gul skjorta som tittar på en stor bit av klippt fisk.
Unga kvinnor mediterar i skogen, bär arbetskläder och en cykelhjälm.
En kran som flyger precis ovanför en vattenförekomst
Mannen i halmhatten röker en cigarett.
En ung pojke i en blå jacka svänger ett slagträ mot en boll.
En man som tittar på råvaror.
En pojke i grön och blå skjorta sitter inne i en jordgrävare.
Stor brun hund hoppar över en mindre svart hund.
En gul lastbil med Casterol branding leder en vit lastbil och blå lastbil ner på vägen.
En publik tittar på början av en drag race vid skymningen.
En person som bär clownmask kliar sig i hakan.
Flera personer lagar mat vid en grill i ett kök.
En äldre asiatisk man tittar på en kamera i en stor samling människor.
Folk jublar som en cyklist rider sin cykel från en ramp
En man rider en mountainbike på en skogsstig.
En polis står och patrullerar i hörnet nära en röd brandpost.
En person som bär hjälm börjar åka skateboard nerför en gatukulle.
En person går i en stad med en grupp fåglar.
Två barn leker i en hög med ospolat toalettpapper.
En tjej i svart klänning och orange jacka.
En arbetare sopar vägen när en maskin kör framför honom.
En man hoppar in i en inskärmad utomhuspool.
En målvakt dyker för att förhindra bollen från att gå in i målet.
En svart hund i vattnet.
En man med vit hatt, vit skjorta och svart förkläde grillar kött.
En flicka som sjunger och dansar med en rosa hatt på.
Tre barn alla bär capri byxor och långärmad huva jackor ivrigt väntar på ett tåg.
En stor grupp av cyklar racing på gatan
Män och kvinnor i baddräkter sitter utanför en stock svett lodge med träd i bakgrunden.
En man som sitter på en bussbänk och lyssnar på musik.
En brun hund sniffar en vit hund framför två kvinnor.
Folk spelar i fontänen en solig dag.
En cyklist som gör en somersault med cykeln framför en publik.
En man som hoppar från en byggnad till en annan i närheten
En skulptör flisar bort i marmor för att skapa en staty.
En man och en kvinna går in i en buss och betalar vägtull.
Det finns en dam som bär hennes resväska bakom henne på vägen.
En man i mörk skjorta och glasögon håller en mikrofon.
Fyra personer åker rullskridskor med åskådare i bakgrunden.
Den orangea ryttaren kör en motorcykel på ett hjul.
En brunettkvinna med mörka glasögon och en röd blus äter.
Två hus och eld
Två flickor i röda fotboll uniformer som springer efter en fotboll.
Två skateboardmän i hög hastighet.
En svart person i svart och rött sover på en bänk med ett öppet svart paraply.
En kvinna i blå kostym vänder sig till andra i ett arkivrum.
En man håller i en gitarr med ett ljus som skiner bakom sig.
Stor vit hund som springer på gräs
En brun hund springer genom vatten och bär en boll i munnen.
En svart och vit hund hoppar genom vattnet.
En flicka i rosa klänning står på huvudet.
En man utför ett skateboard trick.
En man går in på en transportstation och två officerare i neonjackor står vakt.
En liten flicka som rider på en gul leksaksbil i plast.
En ung man hoppar upp från sin skateboard på gatan framför ett hus.
En äldre kvinna arbetar i ett eftergiftsstånd.
En ung pojke hänger huvudet ner i ett däck sving med grus under.
Flicka som cyklar på en gata nära många butiker.
En ung dam i randig skjorta väntar på den unga damen med blont hår som skriver.
Kvinnor som spelar volleyboll i sanden nära havet.
Kvinna med grön skjorta och blå väska stående på en trottoar.
En man med hatt inspekterar en annan mans tatuerade arm.
Två dobermaner slåss eller leker tillsammans på en gräsmatta.
Två män hängande runt en byggarbetsplats.
Två män som arbetar med trä på ett jordgolv.
Orange hund går i grunt vatten.
En kvinna som hjälper en liten flicka att välja ut och läsa en bok.
En ung flicka som bär svarta stövlar håller i staketet och har en klubba.
En hund som simmar längs havet med en bark i munnen.
En pojke skyfflar gödsel i en brand medan en man tittar mot kameran.
En ung kvinna i rosa skjorta som står på trappan ler mot de vackra rosa blommorna.
Kyrkomedlemmar ser en pastor hålla en predikan.
En fotbollsspelare som håller bollen jagas av en annan fotbollsspelare från motståndarlaget
Cheerleaders visar symmetri när de förbereder sig för att utföra.
Cheerleaders i blått uppträder på en fotbollsplan under en gul fotbollsmål stolpe.
Cheerleaders bär blå promenad på fotbollsplanen.
En man och en flicka tittar båda på något av intresse.
Lokala människor försöker sälja varor gatan sida.
En man i brun klänning som står i sand.
Fyra pojkar leker på en lekplats i trä.
Mannen i den röda overallen står på trottoaren.
En grupp flickor i blå kläder.
En rad cheerleaders i blå kostymer väntar på att uppträda.
En kvinna och ett barn leker på en snötäckt gård.
En hockeyspelare i svartvitt kolliderar med en annan spelare i blått.
Pojke i orange tröja har fotboll och är på väg att tacklas.
En person i blått klättrar upp för en mycket hög klippa, fäst av röda och blå rep.
En man hoppar från en sten i vattnet.
En liten flicka är på väg att hoppa in i en lerpöl med sina blomkängor.
En pojke i shorts sparkar medan han står i grunt vatten.
En stad i centrum där en person lutar sig mot en byggnad medan han använder sin mobiltelefon.
Män spelar ett spel i röda uniformer
En vit hund i koppel bär en gul jacka.
En man på en hiss och en annan på taket av byggnaden tittar.
En svart och brun hund som drar i rött koppel.
Fyra kontorsanställda arbetar med ett projekt.
En stor brun hund och en liten grå hund på en stenig yta med ogräs bakom sig.
En pojke studsar på en studsmatta.
Den svarta och vita hunden föder upp fåren.
En man visar tre barn som sitter vid en bordsskugga.
Tjejen i rosa Hello Kitty-skjorta hoppar.
En motorcyklist lutar sig in i en kurva med sin motorcykel
En kvinna i svart klänning som sköljer ur en trasa i en blå hink.
Två små bruna apor på en vägg som bråkar med varandra.
En person lutar sig på baksidan av en buss, medan två andra människor ligger på gatan.
En ung flicka i rosa sitter på marken.
Ett barn som bär en röd topp står bakom ett blondt huvudbarn som sitter i en skottkärra.
Gamlingen städar trottoaren utanför en affär.
En äldre kvinna med grått hår och glasögon, tar en tupplur i sängen.
En orientalisk kvinna som jobbar på en branschlinje.
En motocross ryttare är på en gruskulle.
Två barn leker på stranden och flickan hoppar.
De två människor som bär grönt sitter ner och omges av tomma platser.
En fotbollsfan som visar sin hängivenhet genom att måla hans ansikte.
En äldre man i blå och vit skjorta spelar saxofon.
Man med hjälm utför ett trick medan rullskridskor.
Tre män, två med skjortor, en utan att arbeta på taket av ett hus.
Två cykelförare står med 3 cyklar parkerade vid bilen.
En man, som bär cowboyklädsel, rider en häst i en rodeo, medan en folkmassa bakom ett barrikaderat staket omger honom.
En man som rider en svartvit tjur medan folk med cowboyhattar tittar på.
Två par omfamnar passionerat på en strand, medan ett äldre par ser på från ovan.
En grupp människor samlas framför ett rött hus.
En ung flicka, i en stjärna och ränder baddräkt, gör en baklänges vända på stranden.
En söt valp hämtar en gul ring tuggleksak på gården.
Folk samlas för att dricka och prata utanför dörren till en byggnad.
En grupp tonåringar spelar musik vid ett utomhusevenemang.
En grupp människor på en rodeo tittar på en cowboy som kastas från en vit häst.
En man rider på en häst när folk tittar på.
Barn, däribland en med ett målat ansikte, klappar små sköldpaddor som kryper i det gröna gräset.
Ett barn med solglasögon och en skjorta fylld med smuts.
En hund jagar en boll som har sjunkit i vattnet.
Fyra barn som leker i vattenpipor.
En kvinna med matchande ljusblå t-shirt och headscarf sitter på en stol gjord av sten.
Ett par beter sig som om de simmar framför en fiskutskärningsdörr.
Två damer i Tutus dansar på gatan.
Ett par kvinnor uppträder på gatan för en massa människor.
Två klättrare sitter på toppen av ett berg fäst vid rep.
Fem personer sitter på hästar på en rodeo.
En vit och svart hund springer på gräset.
En kvinna ler inifrån ett rött tält som är omgivet av snö.
En man med vit mössa och vit tröja som arbetar på ett tak.
Semi-pro kampsporter utövar sina mest kraftfulla rörelser.
Ett litet barn i randiga byxor sträcker sig efter en vit spis i ett rött golvkök.
En cyklist utför ett hopp vid några träd.
En ung man klädd i en jersey och shorts tittar på några Ultimate Frisbee spelare i aktion.
En man på en mobiltelefon med cowboyhatt och en blå och vit skjorta står på en trottoarkant.
En man sitter på en stol, medan många människor går framför honom.
Två små barn hämtar vatten från en stor behållare.
En pojke utför tricks på en tegelvägg med en skateboard.
En man som pratar medan en dam tränar.
En grupp unga damer som går nerför en gata i ett turistområde.
En kvinna spelar ett instrument medan många tittar på henne.
En motorcykelförare vänder motorcykeln på sin sida medan racing.
En äldre man med glasögon i svart jacka och svart hatt.
En ung flicka hoppar i luften framför ett vitt hus.
Stor svart hund och kattunge märkligt tittar på träväv korg.
En ung kvinnlig hejaklacksledare klädd i en blå uniform hejar framför en grupp bandmedlemmar.
Ett band av musiker står på gatan.
En brun hund knaprar i den vita hundens ansikte.
Tre personer på en klippa tittar ut över vattnet nedanför.
En man står och bär lastbyxor, orange hatt och gul skyddsväst.
En man utan tröja spelar tennis.
En man som sitter på en trottoarkant i en park.
En man som försöker slå världsrekordet för att hänga upp och ner.
En kvinna med brun klänning håller ett glas och en cigarett mitt i ett rum fullt av människor.
En grupp byggnadsarbetare går förbi en byggnad under uppförande.
Två byggnadsarbetare, den ena med en gul metallbit, och den andra med verktyg.
En gammal man och hans hund står vid sidan om med en vagn.
Två kvinnor står i sanden i sina bikinis.
Ett barn som sitter i en barnvagn och bär ett stetoskop.
Blond flicka i rosa och vit klänning svänger.
En hund plaskar i en liten pool med en liten fotboll.
En man med mycket smycken och punkrockkläder ställer sig mot en tegelvägg.
Två män lägger armarna och benen åt sidan.
Ett ungt asiatiskt barn äter röd söt bönpasta.
En hund simmar i en pool medan en annan tittar.
Sköterskan är klädd i vitt och går på en gata.
Personens fot vilar på fluffig svart hund.
Äldre kvinna i randig klänning, vit jacka, går nerför gatan med shoppingväskor.
En grupp människor avfyrar en luftraket framför en marina.
En svart och grå hund leker med en blå boll utanför.
En tjej med en gul EL Dorado Elementary School skjorta på att visa storleken på något med hjälp av fingrarna.
En man med paraply sitter på en bänk i ett offentligt område.
Det finns många barn som arbetar med olika aktiviteter i klassrummet.
En pojke i blått cyklar i en skatepark.
En liten flicka jagar en rosa boll över grusuppfarten.
En fotbollsspelare gör en kick.
En grupp backpackers tar en paus under ett närliggande träd.
En trefärgad hund springer på det gröna gräset.
En man som står på sanddyn och sträcker sig mot himlen.
Två barn flinar och kramar varandra.
Person på en skateboard i luften
Kvinna med glasögon som arbetar på en symaskin.
Ung pojke som använder en dammsugare på en matta.
Två röda hundar springer i grönt gräs vid ett staket.
En fotbollsspelare hoppar i sidled i luften för att sparka bollen.
En brun hund som hoppar genom vattnet mot stranden.
En liten pojke omgiven av en hög löv.
Två kvinnor sitter på en soffa med röda och vita kuddar med käppar bredvid dem båda.
En ung blond pojke som ler stående på en trappa
En liten flicka och en pojke klädd i rött äter flingor ur lila skålar.
Två män knäböjer på en trottoar.
Män arbetar med en cementblandare.
En man arbetar på ett stort fordon.
En gammal flintskallig man skriver på ett papper på ett bord.
En man hoppar ner från en sten i vattnet
En ung pojke håller i sig och rider en lina nerför en kulle.
En man klättrar uppför en klippa högt i luften.
En brunett hanunge sitter i ett handfat och håller i en tandborste.
Ett förtjusande litet barn som tittar upp i ljuset.
Två män cyklister undersöker kedjan på en cykel på natten.
Musiker övar som regisserat av en regissör.
En byggnadsarbetare sköter en cementblandare medan han talar på en mobiltelefon.
Arbetare kör en slang bredvid ett hus.
En grupp arbetare utför en del byggnadsarbete.
En man arbetar med elektronisk utrustning.
En man är böjd över att arbeta på ett rött fordon.
Äldre man målar en bild av gamla ruiner i bakgrunden.
En kvinna i kostym och handskar leder en liten orkester i ett ljust rum.
Två vuxna och ett barn väntar på att gå över en gata.
En hund försöker plocka upp ett stort däck med munnen.
Två hundar leker på en åker.
En man i randig skjorta som säljer grönt och gult melon på baksidan av en hämtning.
En grupp unga vuxna på cyklar
En kvinna i svart klänning och höga klackar sätter sig på en cykel.
En person klädd i blått utför en backflip.
En grupp kvinnor har orange bikina toppar och orange saroog kjolar.
Fyra män står bakom kassan och dricksburk.
En gammal man med långt grått skägg sitter på en stolpe med två andra män.
En kvinna som spelar basgitarr på scenen med sitt band.
Den här mannen är fackföreningsanställd och tjänar 95 000 dollar om året.
En man rider en rosaaktig motorcykel på en kulle.
En man klättrar på ett metallstöd i läktarna på en stor arena, vid ett fullsatt idrottsevenemang.
Två personer, en på telefonen, framför ett tåg.
En man pratar på en mobiltelefon bredvid en bil parkerad i en mörk gränd.
Två män med paddlar i vattnet.
En gammal man sitter utanför en öppen dörröppning på en låg pall
Några svarta killar som pratar med en tjej.
En shortspojke står bredvid en vattenstråle.
Två personer slåss i en karate tävling med domare tittar på.
En ung man blockerar en kick under en sparring match, medan domare väntar.
En man som blev slagen under någon form av kampsport tävling.
En person som bär halmhatt och står utanför och arbetar med en stålapparat med en hög kokosnötter på marken.
En asiatisk man i polotröja reparerar en tennissko.
En ung man hoppar med en surfbräda över vågorna.
En svart hund fångar en frisbee i en park.
En svart hund springer på stranden medan en ljusbrun hund hoppar upp för att fånga en pinne.
En smutscyklist landar på en ramp.
En skateboardare flyger över luften medan andra tittar.
En fotbollsspelare bär bollen under en match.
Denna bild visar en grupp soldater i kroppspansar med röda sköldar
Gruppen i traditionella kläder spelar instrument.
En man i randig skjorta tar en bild medan en man cyklar bakom honom.
Tre män arbetar tillsammans för att rengöra ett unikt designat tak.
En kvinna joggar bredvid en hög betongvägg.
Två fotbollsspelare är i kick off position framför en publik.
Ett litet barn med rosa mössa, blå jeans och vit skjorta står på ett gräsfält.
Tre män bankar på metallfat.
Två äldre kvinnor kan ses från en bil som pratar bredvid en vägg.
En man justerar musiken på en ljudblandare.
Hunden till höger stänger tänderna på de andra två hundarna.
Grupp av människor klädda i svart korsning stad gata
En man och en kvinna som går med två kvinnor som sitter i bakgrunden.
En man nickar på ett öra av majs
En kille på Rollerblades som glider över en räls.
En grupp motocross-förare ställde upp för att börja.
Ett fotbollslag i marinblå som springer ut på planen börjar en match.
En ung flicka i svart väst hoppar.
Fans tittar på när spelare vilar mellan sessioner i en fotbollsmatch.
En liten flicka går ut och skrattar.
Det finns en stadion full av människor som tittar på sportevenemang med manliga spelare.
Den perfekta utsikten bakom en fotbollsmålstolpe.
En fotbollsspelare i gul skjorta kastar bollen tillbaka.
Fotbollsspelarna går på planen.
En kvinna sitter baklänges på en stol mitt på ett fält.
Hunden hoppar för att fånga en flygande skiva.
En ung pojke stirrar på vad som verkar vara en gräshoppa när han håller den i sin högra hand vid sitt ben.
Två collegefotbollsspelare står inför rätta.
Det här är damer och en man, i en bar, som delar ut något i en korg.
En sjuksköterska tar hand om en patient.
Två män och en kvinna sitter, armarna vikta, vid ett fönster.
En man som sitter på en soffa och ler.
En servitris uppträder i en restaurang med armarna uträckta och en topp hatt i sin vänstra hand.
En gammal man sitter i en stol och läser en bok.
Två män på ett sjukhus, den ena besöker den andra är en patient.
En man i blå shorts går upp för trapporna.
Tre personer är i ett rum tillsammans och en man har en armsling på sig.
Ett mellanösterländskt par som går nerför gatan.
Skateboardåkaren i den vita t-shirten rider på en träram.
Ett utländskt län med barn på moped.
En kvinna i svart mössa ligger på stranden i en rosa bikini.
De unga männen har trevligt på stranden.
En grupp turister går nerför en asfalterad stig.
En liten flicka på ett rött djungelgym.
En man som bär svarta byxor rider längs en betongkant på rullskridskor.
En liten pojke leker vid en vattenfontän
En blond kvinna i röd topp sitter på en vägg bredvid ett kysspar i jeans.
Motorcykelförare tar en skarp sväng.
En ung man och kvinna i shorts och t-shirts spelar ett videospel.
Fyra kvinnor som dansar på en fest.
Tre byggnadsarbetare sitter runt ett inhägnat område och läser bredvid ett sandslott.
Två personer och en hund som leker i vattnet med en boll.
En man på en vit vattenskidramp på en sjö
En ung kvinna i röd skjorta leker med en kinesisk jojo.
En man ser förvirrad ut när han står framför ett blått och vitt paraply.
En hund springer över marken.
Många lyssnar på en man med mikrofon.
En grupp människor tittar på ett band som uppträder.
Mannen i den gröna jackan framför en sång för en skara människor.
En solnedgångshimle över porlande vatten.
Två byggnadsmän med vita hattar sitter i stolar och läser tidningar.
En man sitter i en vagn med en åsna fäst
En grupp män vilar efter en lång vandring.
En man arbetar under en blå äldre modellbil.
En liten flicka kastar en rosa och gul bit krita.
Två vänner ler och bär stora sombreros.
En man på en stege reparerar bronsbältros på taket i en byggnad.
Fotgängare går runt bilar på en livlig gata.
Surfer gör trick i våg som sett bakifrån
En smutscyklist hoppar genom luften.
En kvinna slår en bit varm metall på ett städ.
Två hundar kissar på brandposten.
Många går på gatan i storstaden.
Skateboarder slipar ett betongräcke.
Tre män i casual klänning sitter på en stenvägg med en till står nära.
Två greyhoundhundar tävlar runt ett spår.
En man i vit skjorta lutar sig mot ett räcke med en kvinna i gul skjorta.
Ett fotbollslag med gröna uniformer och deras tränare kurar.
En äldre pojke dricker ur en vattenfontän medan en yngre pojke tittar.
3 Asiater ritar tecken på papper.
Prarie hundar som ses med, brun svart och vit
En ung flicka går ensam medan hon äter sin väska.
En grupp människor håller tennisracketar, och poserar tillsammans nära ett tennisnät.
Människor med sina ansikten målade för en fest.
En indian i en röd och blå klänning som sitter och plockar på grönt gräs.
Två medelålders män som står utanför ett företag som säljer stolar.
Två personer med vita hjälmar på ridning i en Yamaha röd och svart bil.
Tre killar tittar ut över vattnet med moln i himlen.
Två leende, små barn, ett barn som håller det andra i en gunga.
En person som gör ett språng med sin cykel över en kulle
En man sitter i ett glidflygplanscockpit på landningsbanan.
En man utan skjorta börjar hoppa från en trumma in i en skara andra.
En gammal man i blå skjorta som jobbar på en arbetsbänk.
En mamma tar en bild med sina två små döttrar.
Kvinnan vilar huvudet på handen och sitter i ett trångt område.
En kvinna och en pojke sitter och äter vid ett bord.
En konstnär bär en röd jacka och blå jeans målning på gatan medan han bär hörlurar.
Fyra kajakpaddlare på en moutainbäck.
BMX ryttare bär en svart hjälm får luft från ett hopp.
En kvinna är lite rädd för att en fågel landade på hennes axel medan hon var i lagret.
En pojke skateboardar i en skateboardpark.
Skäggig man i en blå jacka som går nerför gatan.
En gammal man som sover i rullstol utanför en byggnad.
En del människor söker något.
Två unga män som bär potatissäckar drar en dekorerad vagn nerför gatan och tittar på på gatan.
Ett nygift par skrattar under sin mottagning.
En brud och brudgummen dansar med varandra med ryggen vänd mot varandra.
Två hundar leker hårt med varandra inomhus.
En man som ligger på en parkbänk med en flaska alkohol bredvid sig.
En liten flicka i gul klänning går nerför trottoaren.
En flicka som bär gult hoppar över ett rött och grönt rep.
Män i hjälm går nerför en fullsatt gata på natten.
En man i svarta kläder som står på vad som verkar vara ett svart lokomotiv.
En man och en kvinna ler
En brud och en brudgum sitter vid ett träd och ler mot varandra.
En hund som stirrar på slutet av en glasstrut.
Ung man på en trickcykel som hoppar från en murarpyramid.
En kvinna sitter mot en vägg i en tjusig byggnad.
Kvinna i ett fält av högt gräs och vilda blommor som håller upp en gul halsduk
Man paddlar en gul kanot på en flod.
Ung man som sitter på en filt i gräset och äter revben.
En man sågade ett träd och två män plockade upp skräp.
Kirurger observerar en läkare i gröna skrubber utföra en operation.
En man som arbetar med metall och en brinnande eld vid sin sida.
Den här lilla flickan ligger i en hög med löv.
Ett fyra bitars strängband som uppträder.
Mannen i den blå skjortan höll i en kniv och gjorde sig redo att skära i plåtkakan.
Det finns många människor som sitter i grå stolar.
Pojkskridskoåkning på ett räcke på en parkeringsplats.
En del barn sitter på flottar i en sjö.
En man som arbetar hårt på det grova som är gjort av halm.
En cyklist gör ett trick på en ramp.
En kvinna i BH i sängen som sover med ett sovande barn.
Pojkåkning på skateboard, fotograferad från låg vinkel.
En tjej med brunt hår får håret stylat av en dam i en rosa skjorta.
En man tar en dusch.
En man på en motorcykel rider på ett spår och vinkar.
En man som sätter hösnäckor på en kärra.
En brun hund snarkar på den andra hunden medan de båda är i snön.
En far och son njuter av lunch efter en shoppingmorgon.
En liten pojke i badrock sitter på en bänk nära duschen i ett badrum.
En tårtbit serveras på en pappersskylt.
En tjej och en kille mitt i en fältträning.
En asiatisk kvinna som håller ett fan klockor trafiken går förbi.
En man i löpares utrustning knuffar en barnvagn nerför stranden.
En grupp människor sorterar vita och röda väskor.
En man med t-shirt och keps använder en spade.
Pojkar spelar fotboll nära ett mål inlägg.
En hund hoppar i luften bredvid en man på stranden.
En man som står mot en byggnad, i solljuset, som du kan se skuggan av den person som tar hans bild
En man med gitarr i ett band som sjunger in i en mikrofon.
En liten pojke som spelar på gymnastikutrustning.
En kvinna scoopar glass vid ett bord med godis och toppings på den i klara skålar.
En tävlingsbils ljuddämpare brinner.
Kvinnan bär nunnas slöja och äter en smörgås i ett trångt område.
En man i röd uniform hoppar på en idrottsplan
En man håller fast vid något när han dras genom vattnet.
En man gör ett hopp trick på en cykel.
Två män ser på som en tredje sätter tvättmedel i en tvättmaskin.
Folk som spelar, basketboll i luften
Två unga män utför kampsporter framför en basketkorg.
Typ av brud och brudgum skära bröllopstårta.
En indisk kvinna står knä djupt i en vattensamling och tvättar sina kläder.
En grupp människor som såg en stor explosion.
Tre barn väntar vid ett bord på att en kaka ska skivas.
Ett vuxet par njuter av tiden i en bubbelpool.
Flera unga pojkar klädda i orange rock, stående med armarna upp längs sidan en flod med båtar.
Barn drar i ett rep.
Två unga pojkar bär ett stort föremål över ett trädäck.
Vuxna och barn samlades utomhus under ett spräckt tak för att umgås
Barn som bär kostymer sitter framför en iMac-monitor.
En man arbetar med heta metalldelar.
Folk går genom vad som ser ut som ett torrt och härjat fält.
En man som går på en strand som har skräp.
En stor grupp tonåringar mal runt på en uteplats.
Folk tittar på en basebollmatch genom stängslet.
En grupp människor plockar upp skräp på en strand.
En ung pojke springer längs en strandpromenad mot en duva.
En grupp människor, stora som små, på en offentlig plats.
Folk sitter, äter och slappnar av i skuggan.
En sjöman leder en grupp människor medan de är på en båt.
En man med långt brunt hår läser en karta.
Turist som tar en tur bland infödda i den klippiga ravinen.
Man i jeans och tröja hoppa i luften på våt yta som visar reflektion.
En man som hoppar på den hårda marken.
Långhårig man i blå jeans med röd bastrumma ovanför huvudet medan han pratar i telefon.
Rollerblader i grön skjorta och mössa, glider ner för en grön ledstång bredvid stegen
En person som simmar i en swimmingpool.
En man i gul och gul skjorta lägger armen om en man i en blå skjorta.
En man med ryggsäck korsar en livlig gata.
En ensam cyklist som bär hjälm i ett lopp.
PitBull håller en rutig diskhandduk i munnen.
En man som bara är klädd i en handduk ligger i en bastu.
Manlig mc cyklar genom skogen.
Greyhound hund i gul jersey och kör på en grusspår.
En skateboardåkare som hoppar framför en byggnad.
En liten flicka som bär rosa sover i en mans knä när de rider i ett flygplan.
Person i en 3-hjuling som kör på 2 hjul.
En hund som bär nummer fyra springer i ett lopp.
En grupp människor som spelar fotboll bildar en stor hög.
En hona som dricker en skum dryck från en stor, klar mugg.
Någon som har kul på sin surfbräda i det klara blå havet.
En person gör tricks på en cykel i en stad.
Unga flickor som spelar fotboll.
En man med glasögon, en rock och halsduk står framför en blå vägg med en öppen bok.
En kille i blå skjorta sover utomhus.
En liten flicka med blont hår leker utomhus med en liten docka.
En liten svart hund tuggar på fingrarna.
Den ene håller i en öl och den andre tar en bit mat.
Två män och tre barn är på stranden.
En man flyger nerför en trappa på sin skateboard.
En kvinna surfar på internet i sitt hems bekvämlighet.
Två män och en kvinna uppträder på scenen i en "Thomas the Tank Engine" pjäs.
En man i morgonrock står nära ljus.
En leende ung kvinna i orange jacka och jeans, går nerför en vandringsled.
En dam och en man är naturälskare.
En flicka går mot några får i en gräsbevuxen dalgång.
Ett ungt par ligger i sängen.
En medelålders kvinna dammsuger köksgolvet med en behållare.
En häst och ryttare, hoppar en barriär på en kurs.
En brun hund springer mellan två grå stolpar som är mycket nära varandra.
En kvinna med gul axelväska ger en man massage.
En man i en blå jersey kör håller en fotboll
Den vita hunden bär en boll i munnen.
En man som går nerför gatan passerar en tegeldörr.
En smutscykel tar en sväng.
En man med en nummer 12 på bröstet är mitt på vägen medan han kör ett lopp.
En medelålders man som deltar i ett maraton, springer på en gata.
En kvinna i mörkblå hatt och en vindjacka som joggar med hörlurar i öronen.
Tre greyhounds är i en hundkapplöpning på banan.
En dam i blå skjorta tittar på sina tre barn som leker på lekplatsen.
En man utför en back flip medan han förbereder sig för en utomhusföreställning eller tävling.
En brun hund kör över en smuts och gräs bakgrund.
Två tjejer med brunt hår och blå skjortor klappar.
Killen i den vita jackan har en blå hatt på sig.
Fem kvinnor som bär skumma röda och svarta kläder poserar.
Ett gäng löpare grupperade tillsammans med röda och blå ballonger i bakgrunden.
En löpare klädd i rött, vitt och blått springer.
En kvinna i en blå tank topp och spandex shorts springer i ett lopp och en man kommer ikapp henne.
En man och en kvinna, klädd i svartvitt, kör ett maraton.
En man och en kvinna tävlar i ett vägris.
En löpare håller upp ett pekfinger medan hon springer.
En man i svart väst och en kvinna i vit jacka springer i ett lopp.
En kvinnlig vandrare tittar på utsikten över några berg.
En man som följer efter på ett bowlingskott som görs i en gränd.
Två barn som håller varandra i handen och ler.
En kvinna, klädd i gammaldags kläder, syr ett stycke material när hon sitter i en trästol förutom en röd tegelbyggnad.
Minivan kör ner för våta stadsgata på natten, stänker vatten.
En man hoppar från en vårbräda och snurrar i luften med andra idrottare i bakgrunden.
En man som bär jeansjacka ler
Två flickor väntar på gatan medan de bär tajt, knappt där kläder.
En brun hund upp till halsen i vatten
Två kvinnor sitter bredvid varandra vid ett bord i en fullsatt restaurang.
Militär personal med jättesax som står under en "Grand Opening"-skylt.
En kille i grå skjorta och en orange overall som jobbar på järnvägen.
Gamling i svart rock och hatt som sitter mot tegelbyggnad.
En man som står på stranden leker med två hundar.
En dam i jeans och en jacka går bär hennes ryggsäck över axeln.
En folkskara tittar på en helgedom medan de håller sina händer i luften
En man på en rullskoter som håller i repet
Två män som försöker ge vägledning och misslyckas helt och hållet, förvirrar sitt offer i processen.
En grupp människor samlas i ett offentligt område.
En kvinna som bär en svart tank topp och en färgglad kjol tittar på de tillgängliga maskinerna i en tvättomat.
En kvinna på en marknad som sorterar salladen.
En liten flicka med en blå skjorta står bredvid en man som bär solglasögon på stranden.
En man kör motorcykel på ett spår.
En man i blått och svart surfar på en enorm vit våg.
Fyra män som arbetar under en byggnadsställning runt en öppen arbetsplats.
En man i svart skjorta, täckt av paintball smatter, gör ett ansikte.
En surfare vertikalt i en våg med en annan närmar sig honom
En familj leker i en pool och en av pojkarna skjuter något med vatten.
En skrattande kvinna bär en lila fjäderhatt och försiktighetstejp.
Flera människor står på en trottoar nära en man som lutar sig mot en stolpe.
En man jobbar på bygget.
En man som står på betong utanför bär en röd skjorta och grå byxor.
En pojke i röd hatt beundrar en knappt klädd kvinna.
Lång man ducka en tjur i mitten av en arena medan andra människor ser på.
En silhuett av en hund som jagar en annan hund.
En kvinna som svingar tennisracket på en utomhusbana.
Någon använder två stolpar för att vandra på ett berg.
En metallarbetare i en hiss skär en rostig gördel.
En pojke poserar bredvid sin scooter.
Den lilla flickan i rosa äter en burrito.
Karate-klassen ska börja.
En man i blå långa ärmar skjorta och tyg lindad runt huvudet, redo att röka.
En person som utför en kroppslös cykel hoppar över jordramper.
Tre personer är på en vit yta framför ett inhägnat område.
En grupp människor som slutade spela tennis.
Mannen går mot en grupp människor på en lång grusväg.
Två kvinnor som joggar nerför gatan.
De två ljusfärgade hundarna drar på sig ett blått föremål som finns i deras munnar.
En kvinna i blå kjol står när tåget passerar förbi.
Protestanter i en stad som främjar orsaken till att stoppa hunger och krig.
En tackling i en fotbollsmatch.
Kvinnor i lila outfit och man med röd skjorta med hjälp av röd teeter totter
En man i orange skjorta med headset är omgiven av mat.
Två svarta hundar springer i sanden vid en pier.
Två män står på röda sågar.
En vit hund springer i surfingen med munnen öppen
Smutscyklist hoppar nerför kullen.
En boxare med röd hjälm har sprejat vatten i munnen av sin tränare i boxningsringen.
En pojke hoppar från en gunga
Ett barn i randig skjorta sällskapsdjur en vit get som ligger ner.
Den svarta hunden springer på gräset.
En svart hund med röd krage går genom vattnet.
Två män på en crooswalk med en affischtavla bakom sig.
En clown med en röd näsa blåser en bubbla.
En mor sitter med tre barn när de äter glass.
En vindsurfare ramlar av sin båt i havet.
En liten hund som springer mellan gula pålar.
Unge pojke gör ryggsim i en simtävling för sin skola.
En grå hund med mynning.
En individ skrotar botten av sin rätt mat med ett blad de har i handen.
Två unga kvinnor snokar vid sitt restaurangbord.
En vit greyhound hund bär en röd jacka med nummer ett tryckt på den.
En liten pojke i grön tröja som spelar fotboll.
En kvinna sitter på golvet och jobbar på en Apple laptop.
En cykelmekaniker arbetar på att fixa sin cykel innan det stora loppet.
En grupp gymnasieelever går längs trottoaren bredvid en byggnad.
Två asiatiska kvinnor står och pratar vid en gata.
Flera människor rider på rygg och sidor av en bil.
Två män som talar framför en röd askstaty.
Ett asiskt marschband med uniformerade medlemmar i beige, gult och rött spel på gatan.
Flera barn utövar kampsport med trä svärd
En liten flicka är klädd i en rosa ballerinadräkt.
En person är på en ramp på en skateboard.
En asiatisk man med pannband och ansiktsfärg hårt på jobbet.
En man lägger sig ner medan en man och en kvinna tittar åt hans håll.
En kille på en vattenskidbräda gör ett stunt.
En liten flicka som håller i en tennissko.
En ung kvinna med blont hår, klädd i grå klänning, och röda tights, lyssnar på musik när hon går raskt till sin destination.
En kvinna står utanför nära många cyklar.
En gammal asiatisk kvinna sitter framför ett tunnelbanetåg och passagerarna går förbi henne.
En man i luften när han gick ner för en sanddune.
Två blonda hundar står tillsammans på en uteplats.
Små barn leker i gräs nära sprinkler.
En kvinna med en huvtröja och bikini nedredelar som håller en kamera på strandsidan.
Kvinna rider en uppklädd häst på vägen.
Asiatisk polis i blå uniformer står framför en byggarbetsplats.
Lilla scouten lutar sig mot ett fullt utomhusbord med asiatiska matställen.
En man och en kvinna förbereder en måltid.
Två äldre kvinnor som gick över en gata och log.
En vit hund springer genom vattnet till stranden.
En liten tanhund hoppar över ett kedjekopplat stängsel.
Tre hundar är på en inhägnad gård och en hoppar från stängslet.
En blond kvinna som går en plaza framför färgglada byggnader.
En fotbollsdeltagare försöker slå en boll medan en motståndande lagmedlem springer bakom honom.
En flicka med rosa hår borstar sig själv.
En man sätter på några arbetshandskar när folk sätter upp bord för en händelse.
En motorcyklist som gör ett trick i luften.
En blondhårig tjej sätter på sig en cykelhjälm med ett klistermärke som lyder "cool katt" som visas på den.
Person som cyklar på grusspår i skogsområde
Många fotbollsspelare springer på gräsfältet.
En fotbollsspelare som fångar fotbollen.
En fotbollsspelare försöker få bollen från en annan fotbollsspelare som kör.
En asiatisk kvinna spelar trummor.
En man i svart t-shirt och blå jeans drar sig upp med armarna på en stor järnstruktur.
En man försöker fånga en baseball.
En man på en cykel bär hjälm, logotypskjorta och pekar på dig.
En ung pojke leker i vattnet vid havet.
En vit kvinna i vita byxor och en svart topp väntar på bussen.
En grupp kvinnor gör en presentation av en staffli.
Tre män gör en musikalisk uppsättning med ledningar och utrustning över hela scenen, och de håller unika gitarr som instrument.
En man i en blå jacka gnuggar pannan.
En man får en kyss från ett litet barn medan han håller ett spädbarn.
Man går nerför en grusväg med affärer på sidan.
Två personer tittar upp från sina mikroskop mitt i en folkmassa.
Tre män har en diskussion bakom en bärgningsbil.
En bil med en kraftigt skadad främre trycks genom korsningen av några personer och en polis.
En affärsman i gul slips ger en frustrerad look.
Tre män, två klädda i gula kostymer, tittar i baksätet på en bil.
Killen med blå skjorta och glasögon, frenetiskt med armar utsträckta kommunicerar.
En affärsman i kostym, verkar vara upprörd, och han nyper i pannan när han sitter inför flera datorskärmar.
Brandmän försöker släcka en löpeld i New Mexico.
Den lilla flickan i vitt studsar på en flerfärgad uppblåsbar.
En dune buggy går nerför en kulle.
En man som bär Astro Boys t-shirt och har baseballhatt städar en pool.
En nyhetsintervju med en man
Tre gruvarbetare på ett fält letar efter guld.
En liten flicka bär hjälm medan hon cyklar.
Två tjejer som rider på en nöjesresa.
En blågrön bil på en grusväg som stänker vatten till vänster.
En man på tunnelbanan håller sina väskor och tittar på en bok.
En man på en motorcykel är silhuetterad av solnedgången.
En man i kockjacka sitter vid ett vitt bord och skriver i en bok.
En orange, vit och svart motorcyklist racing.
En person klättrar uppför en trästege på en mycket brant, taggig klippa.
Hunden hoppar på soffan
En grupp barn sitter bredvid varandra på en grön duk handel material.
En stadsgata visas med fotgängare och en man som står bredvid en matvagn.
Sex män klättrar på en stolpe i vattnet, fyra män är skjortlösa och de andra två bär skjortor, den ena är vit och den ena är blå.
Folk korsar en bro över en vattenförekomst vid solnedgången.
En BMX-cyklist flyger i luften från en ramp.
En man i svart hatt knuffar mot en jättesten.
En man i tröja och blå jeans tar en tupplur på en bänk.
Två unga män tittar på en annan mans skateboard i en skatepark.
En pojke rider en plastsläde nerför en snöig yta.
En grupp skolbarn övar dans.
En man som håller i en vit hjälm springer på en gata.
Två män sopar och plockar upp en gata täckt av skräp.
En medelålders dam med glasögon och en flerfärgad randig skjorta håller ett nyfött barn.
En man leker med en svart och vit hund.
Tjej i blått försöker få en bas löpare nummer 11 ut under softball spel.
En hund hoppar för att fånga en apelsinfrisbee.
En kvinna vid spisen med en blå ugnshandske tar en klunk av sitt vin.
2 Personer med vita hattar tittar över berget
En grupp människor står i sanden och försöker hålla en stor stolpe.
En husky hund som springer genom en gul tunnel på en hinderbana.
Två små flickor leker i fontänerna.
Ett par leker med en liten pojke på stranden.
En ung blond pojke klättrar på en lekplats.
Två vita kaniner är ute på gräset.
Den här flickan är utanför, sparkar löv, på ett fält där det finns träd i bakgrunden.
Fyra unga pojkar klädda i uniform spelar fotboll.
Det finns en kille med hörlurar runt halsen bredvid en kille i en hatt som tittar utanför skärmen.
Fotbollsspelare torkar ansiktet med blå tröja.
En entusiastisk skara människor som sparkar runt en röd boll på ett gräsfält.
Sex ungdomar skrattar och hoppar upp i luften.
Tre män skrattar när en faller till marken med en vit boll.
En person surfar en stor våg.
En brun hund leker med ett vitt fluffigt uppstoppat djur.
Tre bruna hundar på det ojämna gräset.
En man med svart skjorta och vita shorts, tillsammans med tre andra människor, är runt ett pingisbord.
Två fotbollslag spelar ett spel
En blond kvinna läser med en drink i handen och Oreos i närheten.
Två flickor som bär bikins står i sjön.
En ung man gör tricks med sin cykel på en kurs.
Crowd sitter i ett tält efter en måltid.
En äldre person med en tegelvägg i bakgrunden.
En man som gör ett handstånd utanför ett garage.
En kvinna sträcker sig ut ur skottet och lutar sig över halsband och smycken.
En man klättrar uppför berget.
Denna konstnär i res skjorta mejslar bort vid stenen för att skapa ett mästerverk.
Fem personer tittar på något intressant genom ett glas.
En hoppare får en brun häst att hoppa över ett vitt staket.
En person ovanför sin surfbräda på vattnet.
En utsikt från ovan över någon som tar hand om brickor med fisk till salu.
En kvinna som intensivt spelar tennis i en helvit outfit.
En säkerhetsvakt i en blå skjorta som rör sig genom en flygplats.
En man i kostym väntar på tunnelbanan.
En kvinna med rakt brunt hår och en grön tröja tittar på en annan kvinna med uppstoppat hår och stjärnformade örhängen.
Arbetare arbetar för att rensa upp skräp på stranden.
En grupp människor är på ett täckt område talar, och några av dem bär volontär för parker t-shirt.
En svart hund som rullar i det gröna gräset.
En soldats familj går bredvid honom på en stig full av löv.
Människor på stranden med handskar som samlar sopor
Ett par går runt stranden och hämtar sopor.
En kvinna med solglasögon som står vid ett bord med kryddor.
Peeking genom en dörröppning för att se en man som går med en cykel i kvällsljuset.
En arbetare tittar ut från toppen av en byggnad under uppförande.
En mycket stor brun hund leker med en mindre lockigt hårig hund.
En ung pojke i en blå jacka.
En man med hatt dansar runt i ett område fyllt med ljus och graffiti.
De rugbyspelare tävlar om bollen med åskådare i närheten.
Ett par är gift i en kyrka när gästerna tittar på.
En ung pojke som håller i en pumpa mitt i en pumpaplåster.
En lockigt hårad unge kastar yxor på tjurars huvudmålade mål.
Två tjejer på en restaurang äter.
Tre män reagerar som en fotboll flyger över.
En man som tar ett djärvt språng medan han övar sin parkour
En silverbil som körs på en parkeringsplats, medan folkmassor tittar.
En grupp män i etnisk klänning dansar.
Mannen i den blå skjortan kysser en kvinna framför en bröllopstårta.
Tre personer städar upp en strand.
En grupp tonåringar och en grupp vuxna män pratar sinsemellan i ett utomhusområde.
Brunettkvinna som springer tungan över tänderna.
Två vita tjejer håller upp skyltar reklam för en bil tvätt insamling.
En svart bil på gatan bakom trådnät.
Ett barn försöker undvika att ramla av ett får i rodeoringen.
Militär man skakar hand med en man i kostym som åskådare klocka.
En asiatisk man klädd i vit skjorta och blå jeans ger en powerpoint presentation.
En medlem av den amerikanska armén tar emot en utmärkelse från en asiatisk man.
Uniformerade soldater står i kö i en cafeteria och tar emot den mat de har valt.
Man och barn i ett utställningsbås som tittar på något.
En kille sitter på sin cykel med ett hjul i luften.
Två hundar springer på ett fält framför ett hus.
En kvinna och en pojke sitter på en buss.
Tre personer med vita handskar på att plocka upp sopor på en strand.
Två kvinnor ler när de fiskar tillsammans, en med nät och en med fiskespö.
En man i arméuniform som talar med två asiater i kostym.
Flera män av asiatisk härkomst, tillsammans med amerikanska militärmedlemmar, sitter på ett lunchmöte, medan de pratar informellt och beställer sin mat.
En kvinna skakar hand med en amerikansk soldat.
En man i militäruniform pekar som tre andra män tittar på.
Tre soldater i trötthet sitter runt ett bord.
Tre soldater har en diskussion framför en lekplats, medan andra ser på.
Livvakter samlas vid Beach Patrol-stationen.
En person med grått hår och grå utstyrsel ligger ner på en bänk.
Flera personer, somliga som håller parasoller, rider en lång båt nerför en flod.
Två kvinnor och en man på blå och gula platser i kollektivtrafiken.
En ung flicka rider på en häst genom ett spår.
Tre kvinnor som sitter på piren, dricker, plaskar och skrattar.
Tre fotbollsspelare kolliderar i en hast för bollen.
En grupp hockeyspelare glider längs isen under ett spel.
En hund hoppar i luften med en dam som står nära.
En konstnär målar en bild av en kvinna som modellerar med ett japanskt paraply, medan hon står på stranden.
Mannen i den svarta skinnjackan rusar från sin cykel.
Tre kvinnor klättrar upp i ett trådtorn medan de bär små kläder.
Flera människor äter och pratar medan en annan spelar piano.
Asiatisk man som går i en lerig bäck och trycker på ett träverktyg.
Två cowboys på hästar jagar en ung ko med lassos.
En stor byggarbetsplats med många fordon i en stad.
En pojke med gul skjorta och grå byxor som spelar boll ensam.
En grusväg som har träd på ena sidan och kör ner byggnader på den andra.
Två män sitter på en bänk omgiven av växtliv.
En kvinna i rosa byxor som går bredvid en liten pojke som rider på en leksak.
Två spelare rusar under en fotbollsmatch.
En man i orange väst är vänd bort från kameran och reser sig på en buss.
En liten flicka som glider nerför en rutschkana på en lekplats.
En medelålders man rakar skägget i ett rum med vita väggar som inte ser ut som ett badrum.
En medelålders kvinna har somnat på tåget.
Två gula hundar leker i en grön plastpool.
En man dyker ballonger inuti ett bås med hjälp av ett handgjort verktyg.
En ung pojke klädd i slacks och skiktade toppar använder en lövblåsare i ett gräsbevuxen område vid en gata.
Ett barn ligger på marken och gråter.
En liten pojke tittar på saker genom ett mikroskop
En greyhound är aktiv i ett gräsfält.
Liten flicka i en färgstark skjorta tittar på en blomma i ett vardagsrum.
Två små flickor är på en äng och tittar på naturföremål.
Två män klädda i vitt träffade en boll medan en tredje man går upp.
En man ser på när en kvinna städar en pool.
Ung pojke med en liten fotboll.
En grupp människor pratar medan de dricker öl.
Ett barn i röd skjorta sitter mot en vägg med en karta medan man äter.
En liten pojke sover i sin blå barnvagn.
Ett barn rör vid degen på en skärbräda.
En pappa med sitt barn och en äppelpaj.
En man sitter vid ett fönster på ett tåg.
En hund som går genom vattnet vid havet.
En man utför ett skateboardtrick på ett cementmonument i en stadspark.
Två hundar tävlar över banan.
En kvinna sitter och håller i en delvis vävd korg.
Två män på motorcyklar kör på en tom gata.
En man i grön skjorta och svart hatt som spelar gitarr på scenen.
En tonårspojke gör tricks som hoppar över ett räcke.
En gul hund leker med en stor käpp i gräset.
Två paket slädhundar möts.
En flicka står på gatan och viftar med armen när bilar passerar förbi.
En ung man sitter på en stol med en sko av.
En blondhårig kvinna täcker munnen som en man i svart skjorta med händerna.
Tjejen och en pojke som spelar tennis.
Folk tävlar och killen i grått leder.
En man och en kvinna står i en skog.
Två män i svarta skjortor som spelar elektriska instrument i ett rum.
En person som cyklar på en höjd plattform.
En kvinna som sitter på en av de gröna stolarna håller i en mikrofon.
En man och en pojke ser en hund hoppa för att fånga en boll.
En kvinna med lång hästsvans och en man med kort hår njuter av ett skratt medan du äter dessert.
Sitsad gatumusiker i svart derby spelar blåsinstrument utan att någon lyssnar eller tittar.
En man som bär påsar med grönsaker i ena handen och en bricka med grönsaker i den andra.
Vakter på en konsert, kvinna i röd klänning på scenen.
Barnet rider ett fordon längs en gated stig bredvid ett strandområde.
En kille står på sin london turist monter.
Pojken i den röda tröjan kör med fotbollen.
En kvinna som spelar bas.
En löpare i svart passerar en utomhus blomsteraffär.
Unga kvinnor samlas för en liten fest.
Flera personer samlades i ett kök runt en ö och åt.
En snowboardåkare är i luften och gör ett trick.
Många kvinnor i färgstark saris går in i en stenbyggnad.
Två stora brynhundar som ser likadana ut brottas.
En arbetare svetsar lite metall med full skyddsutrustning medan han sitter ner
En cowboy med vit hatt misslyckas med att vred en kalv på en rodeo.
Tre barn leker på strandlinjen med en färja i bakgrunden.
Ett litet barn som hoppar i en hög löv
Två kvinnor och en man står bredvid ett picknickbord täckt av mat och vatten.
Två män skriver i sanden på en stenig strand.
En man ler när han tittar ner på en orange sportbil som står parkerad vid en trottoarkant.
En man i grön skjorta som rotar en kalv på en rodeoarena.
En lejoninna jagar en svart bison över en gräsbevuxen slätt.
En fotbollsspelare springer förbi en tjänsteman som bär en fotboll.
En äldre man, som är pilot på ett plan, ler.
En båt svänger höger i en öppen flod.
En blond person står framför en byggnad med utsträckta armar.
En pojke gör ett skateboard trick.
En ung pojke utför tricks med en skateboard på en skateboardpark.
Män spelar saxafoner utanför en byggnad.
En man gör en skateboard trick, känd som Ollie, över en trappa.
En brun hund är på det gröna gräset.
Två pojkar i blå skjortor som slåss bakom en grå bil och två andra barn.
Tre kvinnor hoppar lyckligt efter att ha avslutat en road race.
En snowboardåkare skjuter upp i luften över vit snö
Två män spelar fotboll på ett gräsfält.
Ett rockband spelar på en Zune scen medan många tittar på.
Ett band som spelar utanför en Zune-byggnad.
Barnen är i parken och väntar på att få prova den stora sprängningen.
Folk klädda som tomten i en klubb med gröna ballonger.
En pojke som rider en Thomas the Tank Motor scooter och en flicka som rider en rosa scooter är på trottoaren.
Löparen har en batman uniform för loppet
En målvakt i en röd uniform sparkar på fotbollen för att skydda målet.
En cykelförare hoppar över en barriär med sin cykel.
En äldre man tittar över en yngre man som svingar en yxa och hugger ved i en fallmiljö.
Två hockeyspelare tävlar på isen.
En liten pojke försöker göra ett hjul.
Surfare på en enorm havsvåg vid solnedgången.
En hund som skakar av sig vatten efter att ha lekt i vattnet med en frisbee.
En liten flicka gungar, en kvinna står bakom henne.
En person i en stor rosa triangelformade kostym vågor som en man och en kvinna klädd i matchande färgglada randiga och polka-doterade kläder leende tillbaka.
En man och kvinna kysser framför en vit staty
En blond tjej i svart cape står med andra barn i kostym.
En man med glasögon och en grön mössa som somnar på tunnelbanan.
Två små vita hundar med munkorg hoppar över ett litet föremål.
En behandlande försäljare står i solen medan andra sitter i skuggan under paraplyer.
En man spelar gitarr och sjunger in i en mikrofon.
Race bilar på natten i regnet.
En grupp människor njuter av en varmluftsballongtur.
Grupp sätter upp för kampsporter kamp.
En surfare rider en stor våg på en blå bräda.
En dam och ett barn i en jordgubbstur
En man i blå skjorta tar en paus från att gräva i en flod.
Tre personer agerar i en pjäs.
En grupp människor med barn uppträder på en scen.
En person i luften på en cykel.
En ensam bergsklättrare som klättrar på en bergvägg
Tyska Shepherd hoppa genom svart båge medan människor titta på
En liten flicka som sitter på en stol spränger en jättegul ballong.
En man som bär en Vegas-skjorta har en öppen resväska bredvid sig.
En arbetare, upphöjd på en utrustning, försöker reparera en stolpe nära ett fönster.
Två unga män hoppar sprudlande på en utomhusplats.
Fyra män med orange västar är på en byggarbetsplats.
Två arbetare går runt en byggarbetsplats.
En man i en tröja med hatt tittar över en bro vid en sjö.
Ett barn drar katten i svansen.
En blond liten pojke med gröna och blå shorts gräver ett hål i våt sand.
Tre hundar leker i gräset nära lekplatsutrustningen.
Kvinnor på fälten som arbetar på en gård som planterar risfrön.
En gammal man ser eftertänksam ut när han stirrar bort från balkongen.
En publik väntar utanför ett tunnelbanetåg, redo att gå ombord.
En person som gör ett cykeltrick över en träramp.
En kvinna i röd klänning står bredvid en flicka som tittar på vatten.
En hund springer över gräset.
En fotbollsspelare viker en fotboll under en match i leran
En grupp människor som bär hattar samlas med stora väskor.
En fotbollsspelare som bär en blå, Samsung sponsrad jersey snubblar över en annan fallande fotbollsspelare bär en röd jersey.
Surfaren är i vågen.
En folkmassa går på en trottoar strax efter det att det har regnat.
En medelålders kvinna i snygga kläder som håller i en kamera.
En man som står utanför framför ett fält med en stor gul säck på axeln.
En kvinna talar in i en bullhorn en kall natt.
Folk väntar i kön för att gå ombord på en dubbeldäckare buss under gatubelysning
En liten pojke leker med sand på stranden.
Pojkar gör skateboard manövrar med en amerikansk flagga i bakgrunden.
En man och kvinna kysser och tar en bild av sig själva.
En man sitter vid ett bord framför en stor väggmålning.
En man som sitter på en tunnelbana.
Flera personer, däribland en ung flicka med rosa topp och shorts, väntar på en busshållplats.
En pojke i grön kortlek springer i sanden.
Ett barn går och han trycker på sin leksak
Pojke och vit hund springer i gräsfält
En kvinna sitter vid ett skrivbord och skriver på en dator.
Två dirt bike ryttare i luften.
Män i ett kluster under ett cykellopp
Den bruna schäferhunden leker med en pinne.
En kvinna som håller i en handväska står vid kanten av en klippavsats och tittar ut över träden.
Ett par som går på stranden tillsammans kommer förmodligen ihåg goda tider.
En kanna och catcher firar slå en annan baseballspelare ute i ett proffsspel.
Fem personer sitter runt ett bord och tittar på några papper.
En stor skara människor, somliga med händerna i luften, samlas i en stor byggnad.
De fem personerna står under tre solbrända valvbågar.
Två kvinnor kramas medan en tredjedel kliver ur bilen.
Tre kinesiska kvinnor diskuterar något.
Två kvinnor går över en bro över en smal vattenväg.
En man klädd som en clown som cyklar i ett lopp.
En liten pojke i overall glider nerför en orange rutschkana
Många människor njuter av en konsert.
En grupp människor står längs en mur och väntar på något.
En man håller upp handen med en flagga.
Ett barn staplar glatt sina legos nära sin spelplats.
Den vita ankan simmar med en svart hund
Militären arresterar en man mitt på gatan.
En man som samlar halm för att göra hyddor.
Två kvinnor med hattar och en man som knuffade en barnvagn passerade en spabehandlingsanläggning.
En man som cyklar på en offentlig bänk.
En man hoppar en sten på en orange dirt bike.
Tre musiker sitter på stolar och spelar sina respektive instrument.
En liten pojke i en blå huva snurrar handtaget på en vevdriven maskin.
Tennisspelare ses samtala på banan.
En tjej klädd i halloweendräkt bär godis och en lie med en jack-o-lykta på någons veranda i bakgrunden.
En man i flanellskjorta skär en sten.
Ett barn klädd i lila och en vuxen klädd i svart.
En tjej som gör en kick nära en kvinna.
En medelålders blond kvinna riktar ett föremål mot en vagn.
En snowboardåkare som maler ner en sidoskena.
En ung pojke med blont hår leende medan poserar på en trädgren.
Fem pojkar som leker ute på en inhägnad bakgård.
Alla är klädda som zombie på den här festen.
Två flickor i röda kostymer leker tillsammans.
En man i en polisdräkt bredvid en man i en zombiedräkt.
Män och kvinnor i halloweenkostym som har ett samtal
En grön dragvagn står parkerad under ett träd i ett skuggat område.
En man på en motorcykel i luften
En grupp medelålders människor med bärbara datorer och bärbara datorer är uppmärksamma på något.
En man som rullade på en metallstång.
Två motståndare manliga spelare jagar bollen i fälthockey.
Två musiker bär på högtalare, gitarrer och musikutrustning.
En grupp amisher står utanför en kyrka.
Man med mask på höjer handen.
En kvinna som badar ett barn i en specialiserad barnbadare.
Två män spelar basket.
En basketspelare letar efter någon att skicka bollen till.
Basketspelaren i blått utmanar spelaren i orange för bollen.
En man i en Ozzy t-shirt tittar på sin frukost med pocherade ägg och rosta med kaffe på sidan.
Två män med kort hår fungerar.
En stor grupp människor protesterar mot något på en gatuhörnare.
Ett par klädda i udda kostymer.
En vit hund med röd krage hoppar upp från gräset.
Två män från motsatta lag som spelar basket.
En man i Miami basket uniform tittar till höger
En vit kvinna som tittar ut genom fönstret mitt på ljusa dagen.
En liten flicka som borstar ett äldre flickhår med en vit borste.
En liten flicka som tittar igenom en tidning.
En man lyfter tunga stenar och staplar dem ovanpå varandra.
Tittar genom en bils vindruta vid en hund som korsar vägen.
En man i rutig skjorta träffar ett träd med en Axe.
En baseballspelare som svingar ett slagträ
En grupp unga män sitter på klippan och tittar i fjärran.
En man som står vid en mikrofon framför en stor publik.
En ung dam som tröstas av en man efter att hon har sett något sorgligt och det har fått henne att gråta.
Man och kvinna står varandra nära medan en annan man tittar.
En kvinna står mitt på en tegelväg.
Ett datorlabb i en skola, fem personer föreställde sig.
En liten pojke som sover på en randig soffa medan han är insvept i en vit filt.
Soldater tvättar kastruller i röda badkar.
En man i orange skjorta och blå hjälm tävlar sin cykel.
Flera ryttare rider förbi varandra med flaggor.
Äldre kvinna i gul jacka, håller skylten säger "DOWN OCH UT" i urbana området.
Mannen med randig skjorta står bredvid sin motorcykel.
En man i blå rock går ett litet vitt djur när en buss passerar i bakgrunden.
Militär personal lär sig att skjuta sina gevär.
Cyklister bär sina cyklar uppför en brant gräsbevuxen kulle.
Medelålders skallig man som sitter och tittar på två datorskärmar.
En flicka i orange skjorta tänder ljus.
Kille och flicka kysser på tågstationen.
En brun hund sitter i lite snö
Två hundar leker med varandra i löven.
Flera personer i ett band hoppar upp och ner till musiken.
Det här bandet spelar på en scen.
Flera människor marscherar och en håller en menorá när han marscherar.
En grupp unga män kastar stenar i ett främmande land.
En pojke som bär en blå våtdräkt rider på en blå surfbräda.
Den stolta hunden återvänder med leksaken den hämtade.
En mycket upptagen stad gata på natten med cyklister och taxi på vägen.
En man med blå sportjacka och en annan med grön skjorta tittar mot kameran.
En stor skara människor går i en utomhusmat basar.
En sittande pojke spelar dragspel.
En kvinna äter vad som verkar vara en mussla.
En kvinna med hund går nerför en utomhustrappa, en buss bakom henne.
En beväpnad man som simmar och håller en flaska i poolen.
3 kvinnor lagar mat i ett kök.
En man spelar gul gitarr medan en katt tittar på honom.
Flickor går på gatan en solig dag.
En kock och hans två souskockar lagar en maträtt i en restaurang.
En hund slickar sina läppar i ett rum utan mat i sin maträtt.
Fyra byggnadsarbetare arbetar nattetid i staden vid vattnet.
En pojke och en flicka som dansar.
Flera unga pojkar bär blå hjälmar och blå och röda flytvästar på en flotte
En man får mycket lufttid när han vaknar.
Folk slutför en omröstning medan barnen sitter bakom dem på golvet och tittar.
En kvinna vinkar från två högar torkat majsskal.
En liten flicka leker med en stor, vit pudel på uppfarten bredvid en polisbil.
En hund som jagar en rosa boll.
En äldre kvinna med randig hatt, solglasögon, halsduk och blå rutig skjorta.
En grupp människor som gör upphetsade uttryck med sina händer
En man med rollbesättning använder en videokamera för att spela in en trevlig tillställning.
En ung kvinna bär en "Obama" t-shirt.
En grupp unga kvinnor, en i luften.
Människor som cyklar och handlar sent på kvällen.
En grupp män klädda i kostym står på en scen.
Fyra fotbollsspelare spelar på trottoaren.
Två kvinnor, en som spelar instrument och en som dansar, ligger vid stranden.
En svart man håller upp ett Obama 08-tecken.
En man av afrikansk härkomst bär en grå skjorta och silverring.
Kvinnan sitter på en lång, vit vägg.
Män och kvinnor samlas i en rörig butik, kläder hängande på rack är utspridda i hela
En hund tuggar på en pinne.
En kvinna med halsduk på huvudet går nerför en träpromenad.
Ett litet barn sitter på botten av en rutschkana och ler.
En gammal man tar en tupplur i en rickshaw.
Medelmåttiga, vanliga människor går förbi en anläggning.
Två män sitter på en gräsbevuxen bergssluttning med cykelhjälmar.
Krossande man kikar genom en rad ljusblå och grå uniformerade män.
En närbild av en man som skjuter ett vapen i skogen.
Damen väntar på att städa badrummen.
En kvinna i stövlar sjunger och spelar keyboard från en upphöjd scen till en sittande publik.
En kvinna i klänning som spelar sin akustiska gitarr.
En man pratar på en mobiltelefon medan han håller ett Obama kampanjtecken.
En man som bär en Obama t-shirt och håller i en kaffekopp.
En man i grön skjorta lutar sig i en solstol i ett vardagsrum i ett hus.
En liten racerbil med reklam kör på en regnig bana.
Flera människor plockar genom grödor på en stadsmarknad.
Ett asiatiskt barn bär med sig råvaror i en rund korg nerför den soliga gatan.
En asiatisk kvinna lämnar en taxi mitt i stan på natten.
Folk skriker med sina armar stretchade på natten.
En grupp män och kvinnor är i bröllopskläder.
En liten flicka är extatisk efter att ha öppnat en present på sin födelsedagsfest.
Den svarta hunden springer nerför den gräsbevuxna knollen för att hoppa i vattnet nedanför.
En man och ett barn står i närheten av varandra inom en stamgrupp.
En jägare håller en fågel i ena handen och sin pistol i den andra.
En man i orange skyddsväst som håller upp ett djur han sköt.
Det finns en man som håller i en pistol i ett majsfält.
Fyra män med orange säkerhetsutrustning går genom ett fält.
En ung pojke i röd skjorta klättrar uppför en lekplats klippvägg.
En kvinna sitter och ser en annan kvinna leka i poolen.
En pojke hoppar med en solnedgång i bakgrunden.
Kvinna sms på telefon medan mannen på cykel passerar henne.
En svart man och en stor, gyllene hund är på stranden.
Raftar och en helikopter över vatten.
En människa är i fritt fall från en punkt där andra observerar.
Vid skjutbanan övar en man i grön jacka sin skjutning.
Två män i hustrumisshandlare sitter framför ett gäng döda fåglar.
Barn gör sig aggressivt redo för en fotbollspjäs.
En hund travar med en boll i munnen.
En grupp små barn som leker hopscotch på en trottoar.
Guy klipper gräsmattan och lyssnar på radion samtidigt.
En man i duschen med en mohawk gjord av schampo.
Ett ungt blond barn i vit polotröja använder en tandborste på en grodstaty.
Folk går på en livlig gata.
Ett barn, i en grå huva, med ryggen mot kameran, håller upp en amerikansk flagga.
En ung flicka vandrar bland växter och blommor.
Fyra barn sitter på marken bredvid ett träd som är vitt runt stammen.
Grupp av killar som sitter i en cirkel.
Salyo clownen förbereder sig för att göra en ballong djur för liten flicka i rosa jacka.
Tre män draperar ett rep över en väg.
Två unga män står i ett rum med teknisk utrustning.
En liten fågel sålde något i sin näbb.
En kvinna i blå tröja pekar samtidigt som hon står med en grupp andra kvinnor.
Två män i sviter svänger åt vänster, en håller i en portfölj.
En ATV racer spränger nerför banan och skickar smuts som flyger överallt.
Tre personer går längs en bäck i en djungel.
Två vuxna och två barn cyklar nerför en gata.
Släde hundar drar en släde genom en snöig skog.
En man som bär en gul skjorta hoppar in i en sjö omgiven av två vattenfall.
En pojke tittar in i sitt teleskop i ett gräsfält.
En svart och vit hund på en orange koppel hoppar på ett fält.
En fotbollsdomare pekar på att han leder en fotbollsspelare i blått under en fotbollsmatch.
En man i idrottskläder går över en grön gräsbevuxen idrottsplats medan kameramän tittar på.
Lådor med frukt och grönsaker väntar på en mörk marknad.
En stor grupp människor kör alla Jeeps ner för en två körfältsväg.
Det verkar som om den här mannen förbereder sig för att baka något.
En löpare på väg mot en bas medan basmannen försöker ta ut honom.
Folk i blå kläder bär på förnödenheter.
Här är en bild av afroamerikaner som står med doo-rags på huvudet.
Två personer i bowlinghallen.
En blond tjej med en affisch poserar med en svarthårig tjej.
Tre personer har mycket smink och står tillsammans.
Ett litet barn i en vit tröja gör sig redo att ta tag i stången.
Pojke i hjälm som cyklar i maraton.
En hund springer nerför en fotbit på hösten.
En grupp vänner poserar på en pub.
En flicka sitter på en bänk och håller en uppblåsbar tiger bredvid en annan flicka i en färgglad klädsel.
En kvinna ligger på stranden bredvid sin cykel.
En indisk kvinnlig sömmerska arbetar på ett tygstycke.
En ung man hoppar genom luften från en klippig bergstopp.
Folk flyttar möbler genom andra våningens fönster i en byggnad med hjälp av rep och remskivor.
De tre människorna leker runt med en falsk kniv.
Mannen bär vit hatt och poserar med en blond kvinna och en svarthårig kvinna.
Ett par kramar medan de håller i en plasttiger.
Två barn är klädda som karaktärer i Michael Jacksons "Thriller" video.
Kvinna i solglasögon tillsammans med en man i en safari outfit.
En man i en fin mönsterjacka står utanför en klubb med två damer.
En svart och brun hund som leker i vattnet på en strand.
En flicka i rosa rutig rock går nerför en korridor följt av en annan yngre flicka.
Över huvudet på flera människor som går upp och ner för en trappa.
En man lyssnar på hörlurar som står framför två sönderslitna amerikanska flaggor
Två kvinnor tävlar i ett sportevenemang
Tre skridskoåkare tävlar nerför isbanan.
Barn i badsviten går mot vattnet på stranden.
Två personer går nerför gatan och håller hand på hösten.
En man sitter med sin hund framför en målad vägg.
Grupp klass för kampsport, vissa i uniform och vissa inte, äger rum i en utomhus anläggning.
Unga pojkar ställer upp sig på raden av scrimmage under en fotbollsmatch på en grå dag.
En man fångar en enorm våg på sin surfbräda.
Tre tjejer hoppar på en studsmatta.
En brottare faller på en annan brottare som ligger i en ring.
En sköterska som förbereder sig för att linda in ett nyfött barn.
Person på en cykel som bär en kon hatt, med olika objekt i främre korgen på cykeln och bundna till baksidan av cykeln.
En ung skateboardåkare tittar ut i fjärran.
En grupp på 7 kvinnor och en man i en byggnad som fotograferar och pratar.
En liten pojke som bär en rock begravd upp till sina axlar i löv.
En racerförare ler och ger tummen upp före ett lopp.
En vit man som hoppar i sanden på en strand.
En liten asiatisk flicka med en plastpåse med Musse Pigg inuti.
En man som går nerför gatan.
En svart och vit hund biter på en tallkott på gräset.
En fattig familj lämnar sitt hem med bara några få ägodelar.
Två pojkar leker på väldigt gamla arkitektoniska strukturer.
Män på ett kontor med datorer och en projektorskärm.
En man som bär en t-shirt med hjälp av en dator med en mycket stor bildskärm.
En ung pojke och hans hund låg tillsammans på golvet.
En man som bär en grön skjorta åker skateboard på en ramp bredvid ett vitt staket.
Ett barn som sitter i en lila stol och läser en bok.
En kvinna i ett lopp som vänder ett hörn.
Den svarta hunden som bär en röd krage skakar av sig vatten.
En kvinna i rutig kjol och svart topp spelar en elektrisk fiol.
En man väntar vid sidan av vägen, nära en vattensamling.
En man med glasögon lyssnar på hörlurar och tittar på en datorskärm.
En man dricker vin medan han sitter i en stol.
Ett asiatiskt par kysser utomhus på sin bröllopsdag.
Ett barn leker med färg i köket.
Två barn som leker på sidan av en gammal vit lastbil.
Det finns en tjej som spelar ett dubbelbasinstrument runt andra musiker.
En man i svart kostym, vit skjorta och svart fluga som spelar ett instrument med resten av sin symfoni omkring sig.
En tjej i orange slår bollen i landhockey.
På vattenbrynet finns det barn som leker i ett sprinklersystem.
En liten flicka som bär pyjamas leker med block.
En man kör en röd motorcykel med sin dotter i knät.
En bebis som krälar runt i ett gräsfält.
En ung pojke knuffar en vuxen man i rullstol.
Flera kvinnor spelar musikinstrument hemma hos någon.
En hund plockar upp en pinne med munnen medan han trampar genom vattnet.
Två personer står på en strand och tittar på måsar och surfar.
Två män springer sida vid sida i ett fält.
En grupp människor klädde upp sig och dansade.
Två män och en kvinna sitter vid ett barbord och dricker öl.
Två dykare under vattnet som njuter av sin tid.
En telefonreparatör tittar ner från ovan medan han reparerar sina linjer.
En ung man som surfar.
En pojke i randig skjorta och hatt gör tricks på trappan.
Folk korsar en gata på natten.
En ung kvinna står nära vägen med de röda löven bakom sig.
En man i en klargrön jacka rider en ljusgul motorcykel.
En grupp barn och kvinnor som hukar sig åt sidan en ström av vatten.
En brun hund springer genom en orange tunnel.
En stor brun hund springer längs sidan en svart och vit hund.
En wmoan hoppar från land och ner i ett dike.
En ung kvinna i mörkgrön tennis outfit tjänar bollen.
En person i en röd hatt står tittar på de onrusande vågorna.
En hund springer genom ett fält med en boll i munnen
Fyra små barn sitter på hög pall på en restaurangbar.
En man i svart sjömansuniform och vit hatt spänner ihop händerna och gnisslar tänderna.
En tjej i rosa skjorta som sitter på en röd boll.
En hund står upp mot köksdiskarna och försöker komma in i påsar.
En man och en kvinna som ler mot ett gråtande barn.
Flera personer är i en varmluftsballong poserar för kameran med en flod i bakgrunden.
Folk som sitter på taket och observerar något i fjärran.
En man i en ljusblå polotröja spelar ett arkadspel mitt i en mataffär.
En ung kvinna i en ljusrosa klänning poserar för kameran.
En man i mörk blank kostym spelar piano och sjunger på scen.
Band som spelar inför en publik.
En man i grå skjorta spelar munspel.
Cheerleaders på ett fält övar ett drag.
En ung man i svart jacka som sover på en restaurang.
Person på cykel gör ett trick på vitt fäktning.
En asiatisk kvinna i rosa skjorta och bruna byxor drar på en stolpe medan en liten pojke tittar.
En barfota och skjortlös skateboardåkare rider längs en väg.
En grupp gråhundar tävlar med mynningar som täcker deras näsor.
En man i svart skjorta har en stor buske med grönsaker.
Det finns människor som står och ställer sig bredvid vita tält med sorgliga och oroliga ansikten när de ser sig omkring på brädor och sopor utspridda runt om i området.
Ett barn som bär ett stort föremål på huvudet medan han tittar på kameran.
En man med grå skjorta stämmer sin gitarr.
En man sjunger in i en mikrofon medan andra spelar instrument.
En person som bär en röd halsduk och en svart jacka står framför en liten vägaffär bredvid en motorcykel och vinkar.
Flera surfare rider en våg som närmar sig stranden.
Två unga, leende afrikanska barn i färgglada kläder bär en kanna vatten.
En atelet tar en paus och sitter i gräset dricksvatten.
Isåkare bär blå kostym medan racing mot andra åkare.
En pojke vänder en handknäpp på en gårdsplan.
En pojke i en röd tröja rakar lämnar i en hög.
En man som sitter vid ett skrivbord med en stor hög med papper i knät.
En hund bär en orange väst bedragare lekfullt över gräset.
En kvinna som spelar tennis förbereder sig för att servera bollen.
Clad i galoscher hon balanserar göra snabbt arbete av den uppgift som är nära.
Män och kvinnor går förbi en konstnär på trottoaren.
En man på en blå surfbräda är på en våg.
Två män som håller ut sina armar från sina kroppar.
En svart hund springer förbi ett nätstaket med en blå benformad leksak i munnen.
Detta är en liten blå grön och vit manual.
En man som rider på en brun häst ställer sig framför en bergsscen.
En liten pojke som lyfter handen och står bland en massa apelsinpumpor.
Två personer sitter vid ett bord utanför en byggnad.
Den lilla flickan tacklar en man och gör det universella tecknet för "Touchdown!"
En flicka i färgglada kläder hoppar på en säng med en färgblocksquilt.
Tre Orca valar hoppar i en pool vid Seaworld.
En tonårspojke med en blå och vit uniform som spelar en form av hockey.
En kvinna som håller i en ung pojke glider nerför en vattenrutschbana i en pool.
En grupp killar som håller en annan kille poserar för ett foto framför en släpkärra.
Tre manliga simmare tävlar är ett simmöte.
Ett barn hoppar ner i vattnet bredvid en hög med sjögräs.
En brun hund som hoppar genom gräset.
Den tyska herdehunden jagar en boll.
En schäfer hoppar vänster på patchigt gräs.
Flera människor ler när de bär kronor, klädda hattar och målade ansikten.
En man med röd peruk och andra i kostymer är samlade.
En person i en regnbåge peruk och färgglada kläder visar något för en kvinna.
Gamla kvinna saknade tänder står med metallföremål i handen.
Litet folk står på en havsstrand på kvällen.
Det är fyra elever, en skriver.
Tre flickor sitter vid skrivbord och verkar arbeta intensivt.
En flicka sitter vid ett skrivbord och läser en tidning.
En grupp människor som arbetar i ett UNICEF-lager.
En ung pojke har en grön spade.
En kvinna i gult bär ett barn i vattnet.
Män försöker sälja ballonger och bollar.
En grupp äldre köpmän som säljer spränger ballonger och leksaker längs en gata.
En man som står vid ett mat- och dryckestånd.
En man, en flicka och en flicka klädd som en nunna repeterar i köket framför att göra korvar.
En grupp barn som äter tårta.
Två män, en i svart skjorta och en i randig tröja, kock.
En kvinna med dykutrustning förbereder sig för att hoppa ner i vattnet.
En grupp barn och två vuxna sitter på en bänk.
Två fotbollsspelare sparkar en fotboll.
En kvinna i en maroonsjal sitter och ser ut över ett vitt sken.
Tre tunna kvinnor i färgglada klänningar.
En grupp människor i svarta skjortor som går på våt cement genom en park.
Två hundar leker utanför nära vattnet.
En man som bär vit hjälm är bergsklättring.
En brun hund sitter på stranden.
En liten svart och vit hund tittar på en annan brun hund.
En ung pojke som leker i en pool.
En baseball kanna är bowling bollen.
Cykla ryttare tittar på en olycka med andra sportcykel ryttare.
En lemonadförsäljare i en kontrollerad skjorta sitter bakom sitt lemonadstånd.
En pilot vid fönstret på ett British Airways-plan.
En flicka med armen om en pojke som täcker hans ansikte.
En kvinna som syr på sin veranda.
En man och en pojke brottas inne i ett hus.
De lägre halvorna av två barn som spelar fotboll
En svart och vit hund med en blå hundleksak i munnen går över en gräsbevuxen gård.
En våt bulldog skakar av sig vatten.
Det här är en man och kvinna som håller upp ett äktenskapsintyg.
En vit och svart hund racing på ett spår
Tre barn i blå skjortor som svänger på en gungställning.
Flera barn kikar in i mikroskop medan de övervakas av vuxna.
Två kommandosoldater med pistol vid en trappa och en gammal man med hatt sitter på trappan.
En blond man som hoppar från en klippa ner i lite vatten
En man med röd skjorta och vit smock använder en slaktare smart att skära i en skinnad kyckling.
Två män skojar runt som en kvinna tittar på dem.
En man som bär blå kläder trycker på en båt, som är trä och täckt, med en stolpe, och en kvinna som bär svart är passageraren.
Tre människor skördar gräs från lerigt vatten.
En man är vind som seglar i havet.
En liten hund jagar en annan över gräset.
En snowboardåkare flyger från ett hopp som ligger bredvid ett stort rött atomtecken.
Diners sitter vid borden i en restaurang.
En äldre man i brun kostym vilar på en bänk vid vattnet.
Två bruna och vita hundar springer över gräset.
En man med gröna hopp med skateboard på gatan.
En liten flicka som sitter på en plats.
En ung flicka tittar in i kameran, när en grupp människor, möjligen en familj, samlas på en bakgård.
En ung brunett man hoppar över ett metallräcke medan han ler.
En suddig bild av en man i grön skjorta och bruna byxor.
En man går längs sidan en gul cykel på en trottoar.
En man i en blå tröja pratar med en gråhårig kvinna.
En man som kör motorcykel längs trottoaren.
En brun hund som hoppar ner från en sten i en sjö.
En medelålders man tittar på den medelålders kvinnan.
Tre unga pojkar, en ung flicka och en liten hund leker i ett fort av pinnar.
Folk går nerför en ramp i en underjordisk tunnel.
En surfare rider de kraschande vågorna medan en annan följer efter.
En man ligger på marken och fixar ett däck.
Man rider en mountainbike gör ett hopp i luften.
Små tysta vita hundar springer i gräset.
En kvinna med blått ansikte vilar fingret bredvid näsan.
En hund springer genom skogen.
En grupp människor står på en veranda, och en av dem klappar en gul hund.
En ung man som står i ett trångt område.
Tre pojkar i matchande bågar och västar som uppträder med en grupp.
Två kvinnor kysser kinder medan de håller i blommor.
Två vackra damer visar upp de låga snitten i sina klänningar
En flicka hoppar in i en hög med löv
En man i glasögon, en blå skjorta med svart jacka och ett leende
Två män poserar för en bild på en kameratelefon.
Två män med solglasögon på huvudet vända mot varandra i en folkmassa.
Högskolestudenter som sitter på golvet och hejar på något.
En kvinna klädd i en röd tröja, klädd i ett vitt förkläde, och tvätta en stor kastrull i ett handfat.
Blurry människor går i staden på natten.
Två män arbetar i ett kök och lagar pizza i ugnen bakom dem.
En äldre man sitter på en bänk vid busshållplatsen.
En äldre person med vit hatt läser en tidningsbok.
En dirt bikeer är luftburen framför en publik.
En äldre man i rosa skjorta och svart väst spelar flöjt när han tittar på sin not.
En grupp motorcyklister i ett lopp.
En man med gul skyddsväst hjälper till att förbereda ett flygplan.
En samling människor med datorer och videokameror.
Två vuxna i hjälmar leker runt med bergig terräng i bakgrunden.
Två bruna hundar på ett gräsfält, en som hoppar för en boll.
En man som läser ett papper bredvid lagrat fläsk.
En hund går över en vattenpöl i Las Vegas.
En kvinna i röd och svart jacka och en cykelhjälm sitter på en mountainbike.
Fyra kvinnor står tillsammans och poserar för en bild.
Mot en panoramabakgrund från en bergsvy fotograferas en kvinna med cykelhjälm och solglasögon.
En person i grönt surfar en våg.
Två personer är i ett tält nära en tegelvägg.
En man vid sitt skrivbord läser från sin datormonitor.
En kille klädd i rosa och en kille klädd i svart sitter och pratar, en av dem dricker något.
En man som kör en vagn och säljer godis av något slag.
Tre män står på en klippa med utsikt över bergen och havet.
En man i svart hatt tittar på bilder med en annan man.
En kvinna, i randig skjorta, håller på att bada ett barn.
En man i vit rock står och pratar med människor som sitter.
En man i brun skjorta och jeans gör ett trick på sin cykel.
En kvinnlig gymnast i svart och rött tränas på bar färdigheter.
En man i mestadels läderkläder står i ett nöjesområde nattetid.
En man och två kvinnor klädda i vampyrdräkter
En man i röd skjorta sitter på toppen av ett stenigt berg.
En liten pojke med regnstövlar tar en promenad i parken.
En kvinna som håller upp ett barn och gör ett roligt ansikte
En man försöker knuffa en annan som bär en boll.
Två unga flickor, en i svart och en i blått, övar på balansbalkar.
Fem kvinnor och tre hundar poserar för en bild.
En man med en gul skjorta och guldsolmask i ansiktet.
Två personer klädda som djur poserar för kameran.
Barn i en grå huva som står på botten av en röd plastslide.
En person som vinkar hänger på en lina.
En dam med glasögon håller ett barn som tittar upp på henne.
En liten skara människor som hoppar upp i luften.
En kvinna med rosa smällar och ett barn sitter vid ett bord, på väg att äta en måltid.
En man med gul skjorta sjunger in i en mikrofon.
En mörk hy man i gul och maroon skjorta fungerar kontroller av en maskin.
En hund står på en cementplattform och tittar ner på spillror.
En hockeyspelare försöker göra ett mål medan målvakten och en annan spelare tittar på.
En vit hund som springer i fallna löv.
En mörk brynhund håller en orange boll i munnen medan han går genom vattnet.
En man hjälper en annan man att vända ryggen på en gård.
Två personer i två kajaker paddlar på kusten, med träd på en kulle i bakgrunden.
En man i en brun trenchcoat som pratar med en säkerhetsofficer i ett köpcenter.
En man med brunt hår med glasögon på att titta upp på någon och skratta.
Fem personer inspekterar cyklar utanför ett skogsområde.
Mannen bär en röd, svart och vit jacka ridandes en cykel nerför en asfalterad stig i en park.
En ung pojke leker i löv.
En man håller en mikrofon i munnen, bakgrundsbelyst av grönt ljus.
En konstnär arbetar på en staty.
Markbaserade militära styrkor förbereder sig för att ge sig av på natten.
En dam med rött hår lagar mat.
En man glider på en betongbänk på sin snowboard när folk tittar på
Folk handlar på en asiatisk marknad.
En person i rött ligger på en bänk i en park, och två par sitter på andra bänkar tillsammans.
En man kajaker i grov vatten.
En man i en blå tröja sparkar en boll medan en annan man tittar.
Ett olyckligt litet barn som sitter på trottoaren.
En man som bär jeans arbetar för att göra en skulptur i sanden.
Rugby spelare tävlar i en match.
En man simmar i poolen med ett barn i flytväst.
Dessa två barn och hundar springer genom ett fält av gräs.
Fiskmåsar överger sin klippa när en våg störtar mot den.
Det är många på berg-och dalbanan.
Ett litet barn som balanserar en tallrik i luften på ena armen.
Två kvinnor står nära en vägg full av annonser.
En brudgum som håller upp sin bruds tåg för att se till att det inte blir blött på en regnig dag.
En bröllopsfest ser på när bruden och brudgummen kysser varandra.
Ung kvinna i sommarkläder hoppar upp och ner på stenig strandlinje.
Ett lag roddare roddar i en grön och röd båt
En man i en skjorta med blommor tittar ner.
Två män i blå overaller, en med bandage.
En kille i marinblå och gula shorts hoppar in i en pool.
En grupp på fem unga vuxna som ligger inomhus.
En monsterbil svävar upp i luften på en arena.
En liten flicka bär hjälm och förbereder sig för att åka skoter.
En grupp barn leker i en vattenfontän.
Ett nyligen gift par poserar utanför i sina bröllopskläder.
Ett nygift par dansar med pengar på kläderna.
En godmodig stunt dras på ögonbindel brudgummen, som hans nya fru tittar på, roade.
En brun hund med en svart krage på och hans herre leker runt på sin fritid.
En man klädd i affärskläder står bredvid en orange och grön taxi taxi.
En del människor står, en del går och en cyklar, i en asfalterad gränd.
Två damer och en flicka slumrar under ett skugga träd.
Skidåkaren bär en gul overall och glider över en gul skena.
Basketspelare deltar i ett spel.
Landhockey laget försöker göra mål.
En man ser vågorna från däcket när han knyter ett rep.
Ett tungset par som sitter i gräsmattan stolar på gräset med en brun hund vid sina fötter.
En fäktningskurs äger rum på en basketplan.
Skaterpojken gör ett trick och får sin bild tagen i luften.
Två män som spelar hockey på isen.
En man som ser på som en kvinna i en brun rock pratar med en annan kvinna i en grå rock.
Tre flickor står tillsammans och gör fredstecken med händerna.
Barnen leker med löv på hösten.
Pojken hoppar upp i luften.
En ung pojke som bär en blå och röd jacka räfsar löv.
En hög med stenar och en grupp människor runt det.
Person som gör ett trick på en skateboard i en skatepark medan folk tittar.
En man och kvinna dricker öl utomhus på natten.
Fyra infödda barn uppträder för en grupp människor.
Någon tar en brun kanot ner till sjön.
Ett par har utsikt över ett torg vid solnedgången.
En man och en varg i arktisk snö.
Två unga flickor som skrattar på en däcksväng.
Manlig gymnast på ringarna.
Ambulansen på lastbilen var i en kollision.
Tre kvinnor sitter på en grön bänk och tittar ut över kusten.
En tjej i röda byxor som rider på en moped.
Fartygsarbetare poserar för en bild i flytvästar på gång.
En man njuter av en karneval spel medan hans vän ser på.
En person leder tre hästar bort mot solnedgången.
En närbild till en stor unik typ plan med en ensam kvinna i centrum.
En man bär en t-shirt som visar en bebis som sätter på en uppstoppad björn.
En cyklist försöker sig på ett trick nerför en trappa utomhus.
En publik samlas runt en man som tittar på en föreställning.
En liten flicka i blått ler medan hon spelar på en repsving.
Ett barn och en vuxen som tittar på varandra.
En kille med svart skjorta och jeans, sittande på en soffa, med flerfärgade fjärilar på väggen bakom sig.
En indisk dam vid en väv som gör en filt.
En skara människor står framför italienska stil byggnader.
En hund fastkedjad vid en stol med skjorta och hatt på.
En person som bär en röd skjorta faller från en vit surfbräda.
En kvinna klädd i grått, sittande på ett picknickbord vid en barnvagn.
En kvinna i en grön tank topp rider ner för en festival rutschkana.
Tre barn står framför två stora däck.
En ung pojke sitter på en skateboard mitt på gatan.
Barn som spelar ett informellt hockeyspel
Ett barn som bär en blå skjorta går på gatan och håller upp två fingrar.
Två personer surfar efter kläder i en butik.
En butik är stängd och en tjej kikar igenom den och tittar på underkläder.
En kvinna i röd klänning pratar på en mobiltelefon.
Två personer med cyklar, en framför löpning med cykel och en i back ridning.
Koka varma paprika på den kalla vintern!
Två motorcyklister rider solbränna på en biek längre ner på gatan.
Unge i blå skjorta gör ett trick på sina rullskridskor.
En skara människor samlas i många olika tält, av vilka de flesta har vita tak, utanför.
En grupp människor roddar en båt i en tävling.
En grupp gamla män som går nerför gatan
En man visar en stor hammare.
En ung mörkhyad pojke i en stor skjorta som sitter bredvid en stor hög med sandaler.
Flera pojkar klädda i mörka färger sitter ner.
Två små barn, en pojke och en flicka, går nerför en trägång genom skogen.
En pojke på gatan har en låda.
En dam i röd tröja och en blå jeans kjol bowling med en orange boll.
En grupp människor rode sig i en båt nära en stad.
En liten pojke i en pool ger tummen upp till kameran när en annan simmar iväg.
En skateboardare är i luften mitt i ett trick.
Mannen svänger med vågen på sin surfbräda.
En officer som slår en man till marken när andra flyr.
En man i blå kläder bestämmer sig för att ta sina privata områden mitt i en protest.
En ung pojke sparkar på hösten löv under fötterna.
En man i solbränna är en av de personer som sträcker sig ut för att fotografera paraden, som har lämpliga män med portföljer.
En ung flicka sitter på en bänk nära ett träd och polerar en sko.
En svart hund med röd krage sniffar marken.
En pojke som spelar hockey ligger på isen, skadad.
Folk får mat från ett matstånd vid vattnet.
En svart man sitter på en restaurang.
En ung flicka sparkar en fotboll i gräset.
En hund springer med en stor tallrik i munnen.
Två män sitter på bänkar och tre män står upp.
En cricket fladdermöss har bowlats ut mitt i stubben.
Kvinnor klädda i korta kjolar ska på fest.
Två collegekillar som lagar mat i köket.
Fyra barn står utanför i en kö i en krabba position.
Fotgängare och cyklister som korsar en livlig gata
En lycklig familj sitter runt i en cirkel i sitt vardagsrum leker med en uppsättning dominoes.
En ung man som parasailerar i havet.
En afrikansk pojke i traditionella kläder tillsammans med två andra pojkar och en kvinna
En motorcykel som slår en wheelie framför en grupp människor.
En basketspelare i vit uniform gör ett hoppskott mot ett lag som bär svarta uniformer.
Tre små flickor ligger på vita kuddar.
En kvinna i lila topp går en cykel mellan två stenpelare.
En svart och vit hund som simmar i poolen
Flickan som bär den rosa randiga skjortan står i dörren med armen utsträckt.
Det finns tre vandrare i närheten av ett berg.
Sex hundar tävlar i en tävling.
En man svetsar något på ett brännblock.
Marinsoldater står längs en röd matta och hälsar på när deras överordnade går förbi.
En hejarklackstrupp som uppträder inför en publik
En gammal kvinna i en lång vit kjol går ut ur en affär på en stenväg.
En hund springer genom ett fält.
Tre personer klädda i rött och svart står på en trottoar framför en beige vägg prydd med graffiti.
En brun och svart hund som simmar i en flod
En man står vid strandkanten på stranden med 4 hundar.
Två varmklädda små barn tittar på ett föremål tillsammans.
Två spelare i rödvit och blå fotboll uniformer huk ner på planen.
Mannen med blå shorts är roddare.
Tre män sitter runt en brand framför en stuga.
En ung pojke rider i en liten båt.
Snowboarder stuntar på sin bräda i snön.
En pojke hukar sig ner, gör en kyss ansikte.
En liten pojke hoppar från en hög med däck i skogen.
En överviktig man som sitter i en lastbilshytt.
Två personer på tunnelbanan sover i hörnet.
Babypojken sover på en filt i gräset.
En surfare som rider på en surfbräda i tuffa hav.
En man som gör ett väpnat handstånd i gräset.
En pojke rider nerför gatan med en yngre pojke bakom sig på samma cykel.
Unga män spelar basket i en tävling.
Två barn dyker sida vid sida i en flod.
En tjej i blå skjorta med en lunchlåda går.
En kvinna är klädd i en dräkt med en stor fjäder i hatten.
Ett par kysser varandra mitt på gatan.
Folk promenerar runt de kinesiska butikssidorna och en man sitter utanför vid ett bord med en laptop och annonser.
Ett tåg går genom en stad.
En man med blå mössa sitter på en pall under ett träd.
Flera unga flickor står på en landsväg.
En man med svarta glas och mustasch pratar.
En bruksarbetare håller på att skala en byggnad.
En surfare i en gul skjorta som rider på en våg på en vit surfbräda
En man bär en röd bandanna
Den tyska herden gräver ett stort hål i sanden.
En liten pojke i blått springer genom en hög med bruna löv.
En pojke på en skateboard är på toppen av en ramp.
En ung pojke som sträcker sig och hoppar.
Folk samlas runt en julgran, bland annat några som bär julmössor, under en julfirande utomhus.
Två hundar springer runt i ett får.
En ung kvinna i en grön tanktopp som går sin hund längs en grusväg.
En mn står på marken, och en står på taket.
Det finns en skara människor i det hektiska hörnet av 18: e St. utanför Bank of America.
Hunden vid stängslet springer på gräset.
En grupp människor tar mat från en salladsbar.
En kvinna som täcker sitt ansikte i skratt vid middagsbordet.
En flicka står på två tunna stockar och fotograferar buffel över en flod.
En man sitter på en upphöjd plattform bakom en dekorativ båge.
Afrikanska amerikanska barn som leker på en gata framför en gul bil.
En man kör med sin cykel.
En grupp ungdomar bygger pepparkakshus.
Arbetare går längs järnvägsspår in i en tunnel.
En kvinna som håller i en väska väntar när passagerartåget passerar förbi.
En liten flicka fnittrar medan hon leker på en leksak.
Två pojkar som äter glass håller en vuxens händer.
Två barn som leker i säckar på golvet.
En basketspelare i en vit jersey förbereder sig för att skicka bollen tillbaka in i spelet.
Någon som kör i sidled på en motorcykel.
En grupp människor som bär olika nyanser av vitt uppträder på ett aktivitetscenter på scenen.
Två unga flickor på lek i ett hem.
Små barn leker inuti ett litet gult och blått rör.
Två småbarn poserar för kameran.
Man i röd jacka ger en tummen upp med ena handen en innehav biljett i andra.
En person viskar till en annan.
Två japanska damer med färgglada kimonor på sig.
En man på en motorcykel tävlar en bil i fjärran.
Två små barn med ullmössor och vantar som täcker munnen medan de viskar till varandra.
En person som gör cykeltrick på en träramp.
En man är på toppen av en klippa med utsikt över skog och sjö.
En man klädd i blått, med en Subway Sandwichskylt på trottoaren.
En hund ligger på sin sida på en trottoar med munnen öppen och visar tänderna.
En äldre man som skär upp ett gäng kokosnötter.
En brun och vit hund har är munnen öppen redo att fånga en grön boll.
En sångare som sjunger med en gitarrist i bakgrunden.
Fotografen håller upp en skiva som har en bild på den som liknar den gentleman han tar en bild av.
En rastamänniska med fasor skär frukt.
En kvinna skriver på en post-it not som är på en tavla full av ljust färgade post-its.
Pojke klädd i röd hatt, blå jacka som skjuter plog i snö.
Två hundar, en vit och en brun, springer längs sidan av varandra nära ett gräsfält.
En restaurang frontlinje, med en varmare fram och en person i en röd Coca Cola skjorta matlagning.
Det finns två motorcyklar med en man och en kvinna på.
En hund leker på stranden.
En blond kvinna som bär förkläde lägger ingredienser i en skål.
En skäggig man och en kvinna i en klänning som håller en kopp.
Två kvinnor med långt hår poserar för en bild
En man och en kvinna ler mot kameran.
Tre män står i en bar med en lila disk.
En man i vit kostym står med två kvinnor.
En man håller fast vid undersidan av en klättring medan han klättrar.
Läkarpersonal i uniform samlas runt ett bord.
En man i våtdräkt surfar på blått vatten.
Arbetare i orange kläder, reparerar en gata.
Två män i orange kläder städar upp sopor som spillts ut på gatan.
Sex grannbarn leker i snön.
Två personer bär näsdukar över sina ansikten, en med blåshorn
En hund står i den vita snön.
Män delar ut mat från en lastbilssäng.
En man i en blå tröja skickar en påse mat till en kvinna i en brun jacka.
Fem män hjälper till med lastningen av en lastbil medan tre kvinnor observerar.
En liten vit fågel tittar på ett litet föremål.
Unga män i vita tröjor, spelar en form av rullshockey.
Kvinnor deltar i en sket på scen.
Två idrottare brottas på golvet i en gymnastiksal när flera andra står nära.
En man i blå skjorta passerar under Samsung båge.
En man under färgglada scenljus spelar gitarr.
En grupp människor vandrar i skogen.
Tre kvinnor och en man har ett vänligt samtal på ett kontor.
En kvinna står på ett podi.
Ett stort antal människor sitter runt flera bord.
Två kvinnor lyfter en påse konserverad mat.
Surfaren gör en vink av en våg.
En man flyger upp i luften med sin surfbräda.
En kvinna som sätter sig vid en vävstol med ett barn som tillverkar tyg.
En pojke och en flicka som dansar med varandra.
Festbesökare på en ravedans vid ett bord med glödpinnar på.
Den blonda kvinnan slår på instrumentet.
En man på nattklubb står i folkskaran med händerna i luften.
Ett ungt par samtalar på en hip dance klubb.
Hundarna springer i vattnet.
Den feta bruna hunden står över den lilla vita hunden.
En kvinna håller sitt barn i ett sjukhusrum.
Flickan simmar är ett blågrönt hav.
Två personer klädda i svarta tröja njuter av atletiska aktiviteter på en övergiven strand.
En liten hund hoppar längs sanden
En man i orange skjorta står vid en krukväxt inne i en byggnad.
En rad människor väntar i elektroniksektionen på en Walmart.
Flera människor lutar sig över sidan av en bro och tittar ner i vattnet.
En man som pratar med en kvinna som skrattar.
Två kvinnor på dansgolvet med andra som dansar.
En kvinna som håller en tallrik vattenmelon på en fest eller sammankomst.
En grupp människor dansar på en mörk nattklubb medan en man spelar trummor.
En man och en kvinna som ler på en nattklubb.
En man i blå baddräkt står på en röd surfbräda på stranden.
En man i brun skjorta och jeans som spelar gitarr och sjunger.
Flera människor klädda i indiska kläder talar med varandra.
Fyra personer går på en strand.
Jockeys tävlar sina hästar på det gröna fältet.
Tre byggarbetare diskuterar hur ett projekt ska startas.
En man och kvinna klädda i gammaldags kläder sitter utanför vid ett bord.
En äldre gentleman åker fast och jobbar framför sitt skrivbord.
En man driver en TV - kamera högt uppe i en fullsatt stadion.
En våt svart hund skakar av sig sig själv.
Man och kvinna bär pälsar medan de går nerför tegelvägen.
En man är på väg att spela gitarr.
En man spelar en grön elgitarr medan han står framför en mikrofon.
3 män i ett band uppträder på en scen.
Två män i svarta kläder poserar för en bild av en färgglad byggnad.
En hund springer över lövtäckt mark.
En person som bär rött cyklar över en grusväg.
En hund med frisbee i snön.
Två män uppträder, en sjunger och båda spelar gitarr.
En skara människor köar utanför en stadion.
Många människor verkar sälja och köpa fisk på en fiskmarknad.
Mannen står bredvid en kvinna klädd som en falsk polis.
En man tar en bild av sig själv och ett skrikande barn i en barnvagn, i en spegel.
Äldre herrar spelar gitarr när de bär vansskor.
En kille med en vit tröja och gitarr drinkar från en burk medan på scenen.
En man som sitter vid ett trumset.
En kvinna i kappa går nerför en trottoar nära Chrismas ljus.
En musiker spelar sin gamla röda gitarr offentligt.
En man i svart skjorta och blå jeans håller i en mikrofon medan ett band uppträder med honom.
En fotograf tar en bild av en fågelmobil.
En hund har sin mun vidöppen försöker bita något.
Två män spelar elgitarrer.
Två män gör handgester och poserar för en bild.
En man spelar musik med trumsetet.
En man går på trottoaren vid en skylt.
Ung flicka i blå klänning och tiara applicera makeup i spegeln.
En kvinna som bär en grön skjorta håller en vit låda framför ett bord med två kaffekoppar nära en annan person.
En ung pojke som håller en pensel över handfatet.
En kvinna skriver på ett papper vid skrivbordet i närheten av betongväggar med graffiti och detritus på ett bord.
Gatuförsäljare säljer olika avdelningar, bland annat ananas och fotbollsbollar.
En man som sjunger in i en mikrofon som en del av sitt band.
Den brunfärgade hunden har en gul leksak i munnen.
Två män skakar hand och ler mot kameran, medan en tredje man står bakom dem.
En man kör en container bredvid några priser staplade i en gränd.
En man och en kvinna går nerför en stadsgränd, flankerad av små företag på vardera sidan.
Två män på kanoter på en sjö.
En stor grupp människor köar och dansar i ett dunkelt rum.
Tre personer står och möter videomaskiner.
Flera män som bär etniska hattar tittar på fotografen på en utomhusmarknad.
En kvinna skrattar medan den andra stirrar på den skrattande.
En polis som bär en gul reflekterande jacka och rider på en motorcykel och viftar med kameran.
En man går förbi en byggnad med många skyltar utanför.
Kvinnor och män protesterar ute på en solig dag med skyltar.
Män klädda i gula jackor ridande motorcyklar.
En man tittar ner på en samling glasblåsta lampor och andra små glasprodukter.
En protest pågår om att rädda våra skolor.
Flera vuxna och barn upplopp för mindre klassstorlekar.
En grupp ungdomar står framför profan graffiti.
En upploppsgrupp bildar en linje bredvid en övervänd bil.
Protester kämpar för barnens rättigheter.
Två unga kvinnor kramar varandra och lutar sig mot en stenmur vid stranden.
Killen i svart och blå våtdräkt surfing
En överviktig man sitter bakom ett rött trumset och leker.
Flickor som spelar basket tävlingsmässigt
En flicka med hästsvans i svart fotboll uniform förbereder sig för att sparka bollen.
Fårhundarna springer i hagen.
En kvinna med röd tanktopp står på en grön matta med händerna uppe.
En man i svart t-shirt och bluesskor spelar bas.
En skjortlös man spelar en röd uppsättning trummor.
En flicka bär en fin klänning och en tiara.
En person simmar i ett grunt turkost hav mot en tom, tjudrad roddbåt.
Protester församlade sig med sina tecken.
En person som bär en svart våtdräkt hoppar högt över en våg med en surfbräda.
Många människor sitter och umgås i grupper på en restaurang.
En racerbil snurrar ut framför åskådare.
Någon gräver i jorden med en spade.
En grupp människor marscherar med pickettecken som hänvisar till skolans budgetar.
Två personer i orangea skjortor hängandes en affischtavla.
En man i svart skjorta och jeans spelar gitarr med slutna ögon.
Två män på en konsertsång.
En kille i en svart huvtröja framför en fabriksskylt pratar in i en mikrofon.
Två tjejer och två män som leker på stranden.
En man klädd som tomten rider i en vagn under en parad.
Folk går upp i rulltrappan.
En kock i en blå skjorta ler framför en stor maträtt medan en medarbetare ser på.
En äldre man står bredvid en kvinna som skrattar.
En man gör hattar av löv.
En konsertmästare som får stående applåder för en stor föreställning.
Två unga flickor med huvudet kikar ut i kameran från en stor hög med löv.
Ett barn bär en röd hatt formad som en hand.
En dam som står i skogen och räfsar löv framför två parkerade bilar.
En man i shorts klättrar upp i ett rockansikte.
En skateboardåkare gör ett högt hopp.
En ung flicka dammsuger medan två pojkar tittar på henne.
En grupp människor samlas i ett rum av en stor rund spegel.
Två hundar tävlar över banan.
Två svartklädda unga män står på trappan framför en byggnad.
Två leende män med sina huvuden vidrörande
3 män i uniform lagar mat på en stor yta.
En grupp fattiga afrikanska barn som sitter i ett klassrum.
En grupp svarta barn i vita skjortor sitter på några bänkar.
Folk som sitter vid ett bord arkiverade med pappersarbete, för en diskussion.
En kvinna i en grön hatt står längst ner i en liten trappa med handväskan i en hand.
En snowboardåkare slipar ner en lång betongskena.
En grupp på mer än 8 talar i mikrofoner.
En snowboardåkare som hoppar från en hög tegelbyggnad.
En man är på scen och sjunger medan bandet spelar bakom honom.
Det finns en orientalisk man som klättrar uppför ett berg.
En man i kostym ser orolig ut när han går på den trånga gatan.
Kören sjunger framför en kyrka.
Fem personer sitter runt ett bord och spelar olika instrument.
Det står en man utanför ett skjul med en primitiv grill som röker.
Två personer sitter på ett utomhuscafé framför en gammal byggnad.
En gammal man i svart trenchcoat står på en marknadsplats.
En äldre dam ligger på en gräsbevuxen kulle framför havet
En grupp demonstranter picket på vägen.
En asiatisk man poserar i en kampsport posera framför en naturlig sjömiljö.
En dam som gör sig redo att knäppa ett foto.
En åsna som bär en massa gräs längs en väg.
En asiatisk kvinna raderar en båt lastad med förnödenheter.
Rader av vuxna som håller en föreläsning i ett klassrum.
En kille surfar på vågorna i havet.
En stor brun hund och en större svart hund som leker tillsammans med en boll.
En man som dricker en dryck och håller en plastpåse långt borta från de andra människorna.
En brottare lyfts från marken av en annan brottare.
En jättelik bidräkt kramar en pojke.
Flickan i rutig hjälper den lilla flickan att mata en häst med ett äpple.
En tjej i baddräkt står framför en randig vägg.
En man i tung rock går uppför en stentrappa med en tung väska med polis i bakgrunden.
En kvinna med vit skjorta hoppar upp i luften och sticker ut tungan.
En man kysser pannan på ett barn som ligger på en soffa.
Vit hund med orange krage promenader på fältet.
En man med stubb i ansiktet håller i ett barn.
Ung, huvad pojke och flicka kurar på trappan utanför stora dörrar.
En arbetare med långt lockigt hår undersöker grönsakerna bredvid broccoli.
En ung flicka som drar i svansen på en alligatorstay
En grupp människor loiterar på en trottoar nära en lyktstolpe.
Man rider på en cykel taxi på en fullsatt gata.
En kvinna i en halmhatt som står framför ett bord täckt av diverse föremål.
Två personer tittar på något i New York.
Folk åker skridskor i en utomhusbana runt en stor julgran.
Kvinna som ligger i gräs med en rugbyboll på huvudet.
Två motocross ryttare sitter på axeln av kapplöpningsbanan.
En färgglad buss stannar i trafiken.
Barn som gick över en hel del av en vuxen till en större byggnad.
Två barn leker i snön.
En man i cowboyhatt kämpar för att förbli på toppen av en beige häst.
Två män står utanför med jackor och kepsar.
En man i blå hatt står bredvid en bil med en spade i snön.
En kvinna i svart går nerför trottoaren.
Flickan klättrar på en konstgjord klättervägg.
Män klädda som tomteklausul går nerför gatan.
En stor grupp människor går uppför ett brant berg med moln hängande i bakgrunden.
Fyra personer med rakade huvuden och vita dräkter som ber.
Ett barn klädd som en elefant som står på en säng som hålls uppe av en kvinna klädd i en Dorothy-dräkt.
Mannen böjd på grå bänk märkt SAN DIEGO, snygg blå soptunna.
Ett barn sitter i en fåtölj i en restaurang och skrattar och kramar Musse Pigg näsa!
En kvinna och ett barn blåser på ett ljus i en muffins.
En man på en gata i tomtedräkt och wrestilng mask.
Ett barn gråter och någon håller fast honom.
Mannen ska ta en bild från det öppna fönstret.
En dam med handskar, och en hästsvans lagar något medan folk står och tittar.
Det finns människor som lagar mat under ett tält och bär stora vita kockhattar.
De två små flickorna hoppar på sängen.
Tre män spelar rugby en av dem bär bollen de är täckta av lera.
Den lilla blonda pojken faller på en säng.
En mörkbrun hund springer bakom en gul hund i gräset.
En lerig hund springer bredvid vatten.
En flock fåglar flyger upp från marken bredvid en byggnad med en väggmålning.
En publik av barn ler och pekar
Två män slåss med låtsassvärd i en medeltida show.
Pojke och flicka bygga metall struktur.
En massa människor på en tågstation.
En dam och en man bär regnponchos.
En liten pojke gråter på en lekplats och lite rider en leksak cykel.
Folk sitter vid ett grönt bord med bordsmattor och gröna glasögon.
Ett mässingsband, med många medlemmar klädda i jultomtens hattar, leds av en man i läderjacka medan man spelar under ett tillfälligt bandskal.
Små barn med händerna i luften
En man i solbränd jacka och blå jeans sitter på en bänk och spelar gitarr, med en annan man i närheten.
En man och en kvinna sitter på stenig utsikt.
Ett par sitter på en blommig soffa medan en äldre kvinna i bakgrunden ler.
En brun hund går ner i grumligt vatten.
En äldre asiatisk man som bär en broderad skidmössa utgör en bild.
En kvinna hukar sig på ett handfat medan hon applicerar mascara.
En man och en ung flicka står tillsammans och tittar på något med ett litet barn i närheten.
Killarna spelar en sport.
Två unga kvinnor klädda i vita skjortor sitter i ett litet utrymme.
Två små barn som blåser bubblor på stoopen.
Den flintskalliga kvinnan står och ler bredvid en rynkande man.
En man och ett barn vid en kassadisk.
Den bruna hunden springer på snön med en vit boll i munnen.
Flera personer samlas runt ett bord i ett lager.
En man hjälper till att knyta ett rött band runt en annan mans högra arm under en gatuparad.
Många samlas inför Lincoln Memorial.
Två personers händer; en av dem gör den andras naglar med en emery board.
En man i hatt spelar xylofon.
En grupp ungdomar som ligger på soffan.
Ungdomar ute på middag på en kinesisk restaurang
Den bruna hunden står i vattnet och skakar av sig.
En man och en kvinna med fjädrar på huvudet dans.
En person på en ATV i sanddyner med en lila himmel.
Två kvinnor knuffar varandra under en rullskridskotävling.
En man i glasögon sitter med huvudet i handen medan han sitter vid ett bord för en asiatisk middag.
En gul bil snurrar bakhjulet medan en man i baksätet tittar.
Människor väntar på ankomsten av ett högt tåg under den kalla vintern.
Två indiska barn som har kul med att berätta hemligheter för varandra.
En kvinna med flätat hår skrattar med en man i röd skjorta.
En svartvit stavordshire terrier har sin tass på stora grenen
Två hundar springer genom ett gräsfält.
Pojkarna och gamlingen delar ved till högen.
En grupp på fem män klädda i solbränna befinner sig mitt i en mycket teknisk miljö.
En man spelar ett instrument bredvid en trummis.
En upplyst matvagn står parkerad på gatan vid skymningen.
En kock tillagar en måltid i ett professionellt kök.
En manlig fotbollsspelare som försöker sparka bollen med höger ben, som den andra spelaren i bakgrunden försöker blockera sin kick.
Ett bobsled team löper genom en snöig stig.
En asiatisk langare med bred konformad hatt med olika frukter och grönsaker till salu.
En gatuförsäljare samlar bröd och kringlor att sälja.
Två unga kvinnor poserar och ler i ett mörkt upplyst område.
En kvinna tar en bild och en annan kvinna står i sidled med armen ut.
En man med mohawk sveper en skatepark.
En man står vid en maskin.
Många människor på en restaurang äter och pratar.
En kvinna tittar över sina varor på en marknadsplats.
Ett litet barn med hatt på ligger på gräset mitt bland några spridda fallna löv.
En liten flicka som tittar in i ett kvinnligt ansikte mitt i en folkmassa.
En man som ramlar av en surfbräda i havet
En kvinna tittar på en tallrik fylld med ånga.
En man och en kvinna vid en måltid, med en hund mellan dem.
Kvinnan i färgstarka kläder dansar.
En liten hund bär en liten kvist i munnen.
En liten pojke leker med höstlöven.
En dam och hennes dotter hoppar i en pool.
Barn som leker i en pool.
Två hundar håller röda bollar i munnen, springer i snön.
En kvinna i rosa håller i en tallrik mat.
Ung person som håller en röd och svart fläkt framför en kampsport klass.
En man använder Wood Silk för att rengöra ett trägolv.
En grupp män i formella kläder talar i en grupp
En kvinna sitter och läser en bok på tunnelbanan.
En hund tar en tupplur mitt i en livlig gränd.
En kvinna äter fisk på en restaurang.
En man och en kvinna poserar för kameran med pungiga läppar.
Mannen filmar ett annat skrivande på en stolpe.
En kvinna som bär en bourgogneärmlös topp och blå shorts klättrar steg till blekmedel
Två rickshaw operatörer väntar på en biljett med trafik i bakgrunden.
En snowboardåkare utför ett stunt i mestadels mörker.
Fyra unga män i ett rum, som arbetar med vissa uppgifter.
En servitör klädd i affärskläder håller upp en stekpanna fylld med kött lastat med sås och dekorerad med citron.
En biker gör ett hopp mittemot en stadsstrand.
En man och en kvinna ler.
Två män tittar mot kameran, medan den i främre pekar pekfingret.
En man utan skjorta står på en scen med eld i bakgrunden.
En man med väst och byxor går över scenen på en konsert.
Den här personen i en vit labbdräkt studerar någon form av genomskinlig scanning.
Två personer går två guldhundar i snön.
Kvinnan hukar sig över en väska fylld med en grön grön grönsak.
Människor och buskar är silhuetterade mot en indigo himmel.
En äldre man som sover i en utomhusstol medan en annan kvinna sitter bredvid honom.
Gammal kvinna med massor av utsmyckade kläder och smycken.
En man rider sin gruscykel genom luften i öknen.
En kille i randig skjorta med gitarr.
En liten pojke och en liten flicka leker utomhus med bubblor.
Tre män står i en skog.
En dam i svart skjorta med rött band och lila kjol på en segerfest
En man i jeans rider en ATV över sand.
En kvinna i röd jacka som håller ett barn i en röd jacka bredvid en cykel.
Två unga kvinnor kramas och poserar tillsammans för en bild.
En liten svart hund med röd krage är i löven med en blå boll.
Nyfödd ligger i sängen något täckt med en filt.
Tre brandmän håller i rep från ovan.
En man som går runt på ett fält och gör vem vet vad.
De två hundarna i snön har ett rött koppel.
Två barn leker med en vit hund.
En liten svart hund jagar en annan liten svart hund genom tjock snö.
En grupp människor är backpacking genom ett gräsfält.
En svart hund och en brun hund som rör vid näsorna i ett gräsfält.
En svartklädd man kör en grön cykel.
En snowboardåkare i klargrön som utför ett hopp på en tävling.
En liten hund som springer på sand.
En asiatisk kvinna står bakom glashyllor med bröd på sig, utanför.
Rådjur och kalkoner står på snötäckt mark.
En blond tjej gillar att äta persika.
Ett barn i röd kortlek njuter av lite konst och hantverk.
Många står på en plattform framför ett tåg.
En pojke med blå vantar gör sig redo att kasta snö.
En liten pojke bär shorts och en jacka drar en röd vagn med en pumpa i.
Tre personer står framför ett skyltfönster och ler.
Man gör en skateboard trick på grön tunna.
En persons hastighetsåkning
En publik väntar på ett tåg när det kommer in på stationen
Ett fotbollslag håller upp en spelare i seger.
En kvinna i grön skjorta och khaki byxor försöker träffa golfbollen i hålet.
Barn på soffan, håller röd duk med vit päls.
En man med tomtedräkt stoppades av två poliser.
Ett litet barn fascineras av en leksakslego i en bokhandel.
En mörkhårig pojke ler medan han ligger bredvid två andra barn.
Ung pojke med blont hår sveper vid bubblor i luften.
En äldre vit kvinna gör muffins i sitt kök.
En pojke är på väg att skicka ner en bowlingboll.
Barnet skyfflar djup vit snö nära huset.
En surfare fångar en stor våg.
Två basketspelare sträcker sig efter en boll.
En man med röd hatt spelar trummor.
En man med en basketboll block ett försök att ta sin boll.
En Miami basketspelare med basket i höger hand på banan.
En man i bara sina underkläder som hoppar på en man omgiven av en massa människor.
En man håller i ett fiskespö och fiskar vid solnedgången.
En man i grön hatt, grön skjorta, bruna byxor och färgglada förkläde vänder en enorm pannkaka.
En man i våtdräkt som surfar.
Två killar är ute på en kall promenad under julsäsongen, kanske för att sjunga.
En ung kvinna och två män dricker öl i en bar.
Medan en bollspelare tittar hjälplöst, hoppar en annan och skjuter bollen mot korgen.
En basketspelare är på väg att lägga sig.
Ett litet barn i säckiga blå byxor springer bort från elden i bakgrunden.
Spelare på en fotbollsplan uppträder för publiken.
Små barn står tillsammans och får ett pris för något.
Två vita hundar med bruna markeringar.
Ett barn i röda och svarta vinterkläder gömmer sig bakom ett snö fort.
En ung flicka med brunt hår spelar schack.
En kvinna tvättar foten i köket bredvid en man i vit skjorta.
En livräddare som sitter på räcket och tittar på vattnet.
En man i lila skjorta med en videokamera på en kvinna som sitter på gatan.
En man som sover på ett plan i ett mörkt foto.
En liten pojke i lila jacka är fastspänd i sin bilstol.
Två pojkar på en båt rider genom vattnet.
En hund som springer med en käpp i snön.
En brun hund som tuggar på en hundgodis.
Fyra barn håller varandra i handen och hoppar ner i en pool.
Fyra barn som håller sig varma under en filt.
En man klädd i tomtedräkt klättrar upp för en stor betongbyggnad.
En svart man med svart hår som skrattar.
En man i solbränna som håller ett spädbarn och en ung flicka sittande på en brun soffa.
En gata fylld med bilar och folk i en stad.
En kvinna som bär plastpåsar går längs en naturskön stig.
En person står vid några trappor i färgglada kläder och glasögon.
Två svarta hundar springer i snö med leksaker i munnen.
En fågel dyker för lite mat.
De två barnen och barnet med den rosa skjortan är omgivna av leksaker.
Matgästerna på en restaurang serveras av en servitör.
En naken man med simglasögon på huvudet med en grupp simmare bakom sig.
Simmare samlas för träning vid en pool med simbanor.
En man i blå skjorta som tar en paus och sitter ner.
Två vita hundar springer med varandra.
En man och två kvinnor som har ett samtal på en gräsmatta.
Människor i vinterhattar står i en tunnelbana tillsammans.
En flicka i en ljusrosa outfit förbereder sig för ett lopp.
Vattenskidare håller linje, mitt-hopp och nästan vände upp och ner.
En man sitter på en soffa och håller ett barn omgivet av barn.
Två kalla människor står nära en stolpe.
En man som säljer varor på gatan.
En man i röd jacka står högst upp på stadiontrappan.
En ung pojke poserar med otroliga hulkhandskar på.
En man klappar händerna med en massa barn som står runt honom.
En tjej i en röd topp håller papperslappar.
Barnet tittar på jultomten.
En surfare gör en sväng på sin bräda.
En kvinna i klänning som gör ett hantverk.
En man och kvinna i masker och kostym skålar inför ett julgransträd.
En flicka hoppar i en pool, med en man som står nära.
En tjej i svart och vitt pannband och rosa slips som håller ett glas med vänner på båda sidor av henne.
En kille och en kvinna med drinkar i handen.
En man och kvinna i svarta rockar är ute medan det snöar.
Ett par klädda i vinterrockar poserar tillsammans.
En man spelar gitarr för ett barn i en sjukhussäng
En kvinna som täcker sig med en handduk dricker en burk vatten.
Tre asiatiska damer går nerför en trottoar med portmonnäer och shoppingväskor.
En kvinna håller ett litet barn i handen och bär påsar.
Två asiatiska kvinnor som sitter vid ett bord och äter asiatisk mat.
Två kvinnor som bär jackor tittar på en bräda.
En person i en tröja sitter och tittar på en bok med ett barn i knät.
Två unga kvinnor som har ett samtal
En stor grupp fotbollsspelare i blå tröjor kör genom fältet.
Två män går framför en grafitti bild av en bil.
Ett barn håller fast sin mor på en släde i snön.
En gammal man och en ung kvinna omfamnar på en soffa.
En person på scen med en ljusshow i rosa och blått.
En korgförsäljare går nerför en livlig stadsgata.
Ett tåg närmar sig i en svagt upplyst tunnelbana.
En pojke i sporttema pyjamas står framför en julgran.
En kvinna i en park står med armen uppe i luften.
Barn är klädda i svarta och vita kostymer.
Flera människor läser vid en lägereld på natten.
En kvinna i grå skjorta som häller en klar dryck i ett glas.
En artist som bär styltor, som är täckta av sina vita byxor, går i en parad.
En ung kvinna som viskar ägg i en glasbägare.
Två unga flickor poserar leende för en bild med en julgran bakom sig.
Tre kvinnor poserar för ett foto framför ett julgran
Två män och två kvinnor håller guldplåtar bakom huvudet.
En spansk kvinna och man i ceremoniell klänning dansar nerför gatan.
En tjej i vit tröja och blå jeans som skriver ett papper på en laptop.
En man glider längs en grön barriär på sin snowboard.
En kvinna med ett tomt uttryck kastar en fotboll som en man i en grå skjorta tittar på sin telefon.
En skidåkare på väg ner för berget.
En svart och vit hund hoppar genom ett fält av brunt gräs.
En kvinna visar sin konst för folk.
Flera människor trängs samman i ett rum med tre stora fans över sig.
Person som gör ett skateboard trick i luften.
Två unga pojkar står i ett kök med trägolv.
Två unga pojkar i kavajer på ett stort fält.
En asiatisk man med en asiatisk unge med en ballong runt huvudet.
En man i röda strumpor som leker med några andra män
Fem flickor i skoluniform går omkring på en platt klippa nära en sjö när en man i bakgrunden sitter på stranden.
En man stoppar i ett lakan på sängen.
En kvinna i rygg och vit klänning som går iväg.
En liten flicka i en orange skjorta med en papperspåse.
En kvinna i jeans förbereder sig för att kasta en bowlingboll i bowlinghallen.
En grupp människor som ska ut och vandra.
Två barn som sitter på en lekmatta och sträcker sig efter något
En gammal man och en bebis i rött.
En skara människor som innehåller en del människor som ler och en del som fotograferar.
En person som ligger på marken under några trappor.
En man i en nissemössa med ett vitt paraply står på trottoaren med två andra män.
Barn leker i snön medan föräldrar tittar på
Två kvinnor som sitter bredvid varandra håller i en bebis och den andra visar sitt armband.
Ett barn som rör vid en kvinnas ansikte.
Ett barn med rosa kläder har en napphållare, och hon sitter på en stol med en annan kvinna.
En kvinna och ett barn väntar med bagage
Två unga flickor klädda i vinterkläder leker i en snöhög.
En kvinna som sitter på en restaurang och pratar på sin mobil.
En orientalisk man med vit skjorta och förkläde lagar mat.
En man fångar en flicka som hoppade i hans armar
Damen har svart rock, handskar och stövlar.
Tre kvinnor poserar för en bild tillsammans.
Den rödhåriga kvinnan i den svarta klänningen har armarna runt en vit man.
Brun och vit hund travning med brunt objekt faller i närheten.
En svart och vit hund med en käpp i munnen simmar.
En flicka håller upp ett gult ballongdjur.
En grupp människor hoppar i luften vid stranden av en sandstrand.
En man och en kvinna som dansar på en scen.
En svart och vit hund springer genom vattnet och håller något rött i munnen.
En kvinna i kappa ligger bredvid en telefonautomat.
Två flickor går förbi ett träd framför en tegelbyggnad.
En man i vit jersey doppar en basketboll.
En kvinna i blå rader en kanot typ båt lastad med växter.
En skara människor sitter utanför på ett torg.
En svart man cyklar tvärs över gatan medan en annan går och håller i en hund.
En kvinna som plockar upp ett barn från golvet
En basketspelare tittar upp och ställer in för att kasta bollen.
En man i hatt och lila förkläde lutande på en metall pizza rack.
En man bär en svart stickad "Paris" hatt och en marinblå skjorta på sidan av gatan.
En man i svart skjorta står bredvid ett tält.
Ett barn i röda shorts som leker i en fontän.
En pojke som äter bredvid ett trähus omgivet av träd.
Två pojkar sitter i en grön kajak på gräset.
En man tänder en stor gnista medan kronan tittar på.
En solbränd hund som springer genom gräset med bakgrunden suddig
En familj i mellanöstern går nerför gatan.
En basketspelare håller bollen under ett spel.
En kvinna som klättrar på en klippa.
Två män som går på en nöjespark den ena trycker på en barnvagn den andra bär på ett uppstoppat djur.
De fyra killarna visas en järnbräda.
En kvinna med röd skjorta läser noter och spelar harpa.
En äldre man tittar ner och ler.
Ett litet barn leker med en liten röd sprinkler.
En man i traditionell klädsel spelar säckpipa.
Två personer i mitten av en smutscykel tävling.
En hund står på en strand vid solnedgången.
De två hundarna springer mot kameran.
En snowboardåkare flyger av ett stort hopp.
En man och en kvinna stirrar på varandra på en balkong inne i en byggnad.
En man i vit sjöman talar med en person som sitter på marken.
En man i en blå kanot navigerar i ett vått land med höga palmfjäder.
En man står på gatan utanför byggnadsställningarna.
Ett lyckligt barn får en hjälpande hand ur lådan med nerf-bollar.
En kvinna i gul skrubb sitter på sjukhus och håller ett sjukt barn.
En hund med en ärm i munnen på en rock som en man bär.
En vit hund som springer på stranden.
Två hundar står i gräset, en springer.
En pojke försöker ta en pinne från en liten brun hund.
Två små barn pratar på ett fält framför en gul varningstejp.
Ung man i en grå tröja som spelar ett gitarrspel.
En grupp på fem kvinnliga barn resonerar utomhus.
Ett barn som bär flytväst i en simbassäng.
En kvinna i svart hoppar i luften på stranden.
Anställda som arbetar med registren i en livsmedelsbutik.
En ung flicka springer barfota på en strand
Tre män i vita rockar tittar på en fjärde man pipa glasyr i kakor.
En kvinna som sitter på en buss med en papperspåse hängande på en bärare
En stadsarbetare som städar sprickorna på en gångväg.
En kvinna, en man och ett litet barn rider en scooter.
Två gamla män har ett samtal.
En liten pojke sitter framför en öppen spis bredvid ett Ginger bröd hus.
Den äldre kvinnan ler när hon håller upp en hammare.
En man, som bär en svart träningsdräkt, hoppar upp i luften och delar sig. På toppen av en bergssluttning visas en stad i bakgrunden.
Två svarta hundar leker hämta med en röd leksak
En snowboardåkare hoppar i bergen.
Den bruna hunden gnager på något i snön.
En kvinna med rött hår som pratar med en gammal man vid vattnet och bredvid en bänk.
En man åker skidor i luften.
En basketspelare som förbereder sig för att skjuta bollen
Miami basketspelare nummer 33 dribblar bollen.
Numret fem Miami spelare dribblar ner i rätten.
Den bruna och vita hunden står upp på bakbenen.
En hund skakar sig torr på stranden bredvid havet.
Snowboarder i luft när du bär gult spetslock.
En snowboard ryttare hoppar högt på sin snowboard i snön.
En hund når för att fånga en boll med munnen.
Tre män spelar basket.
Två kvinnor som skämtar är fångade på kameran.
Ett litet barn ligger hälften på en madrass och hälften på golvet.
Två röda barn låg på golvet.
En kvinna som håller en ung pojke i ett daghem.
En svart och vit hund fångar en frisbee på gården.
Tre personer går på klipporna nära vattnet.
En man i tröja håller i en hammare och ler.
En ensam skidåkare som bär en röd ryggsäck snubblar nerför ett snöigt berg
En man tillbringar tid med sin lille son, som håller i en vit kopp.
En grupp kvinnor delar en måltid i någons hem.
En grupp pf människor och deras husdjur går längs en tågbana
En man cyklar på en grusväg genom svår terräng.
Två män säljer parafernalia som kondomer med Obama-bilder på sig.
En man och en kvinna står i havet och kysser varandra.
En domare stoppar en hockeymatch.
Mannen bär en blå tröja och är barfota på en domstol.
En man med hjälm använder en bankomat.
Två män står vid ett räcke, medan de poserar för en bild.
Tre kvinnor och en man dricker öl vid ett bord.
Två personer springer i sanden vid stranden.
Män som använder spelautomater i kasino atmosfär.
En familj sitter, arbetar och pratar i köket.
Tre hundar leker med en frisbee i snön.
Män i Darth Wader och robotdräkter går på vägen.
En äldre man klädd i kostym står bakom ett guldflätat podi framför en mikrofon.
Ett litet barn springer längs gräset och ler.
Ett rött fordon utanför en byggzon.
Ett barn hålls av en vuxen och sitter på ett bord på ett kafé.
Två hundar springer genom gräset.
En grupp afrikanska barn är klädda i färggranna kläder.
En vit och brun hund springer över gräset.
En kvinnlig skidåkare i en grön med rosa blommor hatt skidåkning.
En fotograf i gul jacka fotograferar en bikiniklädd blond kvinna.
En liten flicka med ryggsäck som sitter ner och tittar på en bok.
En silhuett av en figur fallskärmshoppning vid solnedgången.
Mannen i röd jacka öppnar dörren medan han håller i bilnycklarna.
En hund som ligger på kanten av en vit stol
En skjortlös man är på en blå flotte, som ligger bredvid en gul flotte, som är fylld med last.
En grupp som bär vit poserar för en bild.
En man i våtdräkt surfar upp och över en våg.
En grupp barn som leker i en ström
Två unga flickor leker i ett kök på natten.
Två killar hoppar i luften i ett rum.
En flicka som bär en grön overall och goggles med en vacker solnedgång i bakgrunden
Två kvinnor ligger på golvet och skrattar.
En elefant draperad i rött, blått och guld tyg som går på en stenväg.
En violinist använder en gammal stol som musikstativ
Man i gul tank topp med vän i vit skjorta kolla grillen.
En grupp soldater står tillsammans och bär all sin utrustning.
Ett asiatiskt par har rosenblad kastade på dem av en kvinna.
En grupp människor går genom en skogspark.
En kvinna med kort brunt hår och glasögon skrattar med en brunett man i brun skjorta.
Man med kopp tittar upp medan rider på en rulltrappa
Pojke i grön jacka och en tjej i rött som spelar tv-spel.
En snowboardåkare tar en ramp gjord av snö medan andra tittar.
Fem män som bär turbaner rider på elefanter på en gata i östra delen av staden.
En kvinna står på en vägg för att klappa en elefant.
En grupp kvinnor i röda skjortor som sjunger tillsammans.
En pojke svänger tennisracketen på en tennisboll.
En grupp på fem individer, många av dem barn, stod på en kulle och iakttog ett litet djur.
Två hundar leker hake på ett fält.
Flera personer tar bilder med stativ i snön.
Fem barn på en snötäckt gata.
Den unge pojken slädar nerför kullen i snön.
Det är barn som leker medan vuxna sitter på en bänk.
Två män lagar mat tillsammans i hörnet av gatan.
Fyra byggnadsarbetare arbetar med metallbjälkar.
Det finns fyra snöåkare som går nerför en backe.
En brun hund springer nerför en snötäckt stig.
En vit hund och en svart och vit hund springer genom gräset.
En rullskridskor slipar en räls på en inomhusåkare park.
Två män ser ut som de leker med lådor i ett köpcentrum.
Barn som leker på en lekplats glider nerför en rutschkana.
En grupp på fyra vuxna står tillsammans runt en hög med varor.
En mountainbikecyklist rider på en skogsstig.
En ensam skidåkare njuter av backarna en vacker dag.
En vit hund som går i snön.
Två män klädda i orange dräkter korsar en livlig stadskorsning fylld med bilar, lastbilar och motorfordon.
En arabisk man som går sina tre kameler genom öknen.
En man i brun tröja och en kvinna ler för sin videokamera.
Tre cyklister trampar upp en skogsstig.
En pojke som går omkring på foten av sitt hus och som är gjord av stenar på sina bara fötter.
Två män i blå jackor sitter på en betongstol.
En kvinna i svart våtdräkt surfar i dåligt väder.
Ett litet barn håller i en röd leksakshammare.
En ung pojke leker med leksaksverktyg och bär en namnbricka.
Pojken leker snö.
En liten pojke i khakibyxor som visar en man sin godisröra fylld med godis.
En gyllene retriever går genom gräs med en hundleksak.
En man som bär en djungelhatt vandrar med sin guide i vildmarken.
Ett litet barn arbetar ett färgglatt pussel.
En pojke i grön julpyjamas öppnar sin present.
Flera människor spelar twister vid någon typ av evenemang.
Två barn sitter på en hjortstaty för ett foto.
En pojke hoppar för att fånga en flygande Frisbee.
En blond pojke i ett badkar som häller vatten på sig själv med en gul kopp.
En liten pojke i orange med grå skjorta och khakibyxor som leker i löven.
Ett par och deras barn poserar för en bild framför en julgran.
En liten pojke slog ut flashcards från kartongen de kom in i.
Ett litet barn i randig skjorta som packar upp en present.
En ung pojke i grön pyjamas som leker med en leksak på julafton.
En liten pojke i grön julpyjamas som håller i en låda.
Ett litet barn som leker med sina leksakståg.
Mannen och kvinnan poserar med falska glasögon och mustascher.
Hunden står på något medan snön faller runt honom.
En skateboardare flyger genom luften på en röd skateboard.
En grupp dansare med svart spandex dansar i en studio.
Tre kvinnor sitter på en bänk och pratar.
En kvinna och en man poserar med Groucho Marx förklädnader.
Två kvinnor cyklar nerför en grusväg.
Tre personer är i snön.
En man och en kvinna sitter tillsammans i mörkret, tittar framåt på en stadsvy i fjärran.
En man i sandaler sätter sig ner medan han läser tidningen utanför.
En snowboardåkare i en grön jacka fångar lite luft.
De två männen spelar cricket på en stadion.
Det finns 2 skjortlösa pojkar som hoppar upp från lite vatten och tittar på en fotbollsboll.
En person åker skidor nerför en skogbevuxen kulle.
Brun hund med vitt märke i bröstet och svart krage går över en lem på marken.
Ett litet barn och en hund leker i snön.
En person i en vit hjälm fastspänd i en gul bil
Ett äldre par diskuterar en grönsak.
Man i röd t-shirt poserar med två unga kvinnor och tre ölflaskor.
Tjejer i svarta klänningar som dansar på discot.
Fyra kvinnor står på händerna på ett gymgolv, klädda i samma kläder.
En man hoppar in i surfingen.
En liten pojke sitter på ett steg medan en grill röker i bakgrunden.
Den lilla pojken i den blå skjortan är omgiven av hejaklacksledare.
En man i röd skjorta står med två kvinnor som bär vitt och ler.
Fyra personer poserar för en bild
Flickor, som alla är klädda i klänningar, dansar i ett mörkt rum.
Många människor äter i en fullsatt restaurang.
Någon åker nerför en snöig kulle.
En man som spelar ett spel på sin dator.
En man med vit hatt och brun skjorta, bakom en kvinna i rött, ser åt vänster.
Inne i en bar finns personer med röda skjortor.
Två bruna hundar leker i snön.
En ensam person som står på en klippa och tittar på måsarna.
Två vita hundar leker tillsammans på en något snöig lapp av grönt gräs.
En svart och vit hund springer med munnen öppen.
En kvinna i badrummet i pyjamasen
En pojke som leker i en lerpöl.
Flera olika färgade hundar springer i ett snöigt fält
SMU basketspelare kör till korgen.
En snowboardåkare rider sin bräda från en graffititäckt vägg på natten.
Två personer står och tittar på en ljus skulptur på natten.
En kvinna håller ett nytt barn i gult på ett gammalt foto.
Kvinnan lägger en boll i hundens mun.
Det finns en bild av en grön, vit, svart och röd flagga.
En orientalisk person ro en båt, full av grönsaker, nerför en flod.
En ung flicka som åker skidor nerför ett berg.
Människor på en inomhuskarneval med ett spel med stora fyllda djur som priser.
En man i blått på en arkad spelar ett fiskespel.
Två unga kvinnor surfar på internet i ett café
En person som dansar gör ett danssteg där hela kroppen är på marken förutom en hand.
En grå egret tar en flygtur.
En kvinna som sitter vid ett bord utanför en affär som säger parkering i fönstret.
En slägga får ett ansikte fullt av snö på en sluttning.
Två män sitter i en restaurang medan en av dem håller ett papper upp till kameran.
Tre asiatiska människor spelar musikinstrument.
En grupp på fyra pojkar leker med lera i vattnet och gräset.
Många människor spelar färgglada karneval spel.
Människor står på karneval spel av ballonger och fyllda djur på väggen.
Två personer står utanför en affär på en stadsgata.
Två personer som gör det mellan stenar.
Tonåringar spelar i kundvagnar på ett tak.
En breakdancer visar ett imponerande handstativ i ett kraftigt graffitimärkt rum.
En man i blå skjorta riktar sig till folk.
Mannen är på en skidbåt i vattnet.
En man fångar luft när han snowboardar.
Två ryttare och tre vandrare är på väg nerför en dammig stig.
Flera människor rock vandring med ryggsäckar och promenader pinnar.
En ung pojke i en blå fotbollsuniform som jagar en boll.
En collie hoppar över ett vitt hinder.
Någon är snowboard nerför en kulle, strimlande snö.
Ett barn sitter på ett fallet träd.
En kvinna i brun tröja med några smutsiga skålar i vänster hand.
En pojke bär en grön, blå och grå jacka medan du laddar ett gevär.
En man i blå skjorta kastar en fotboll.
Ett barn håller upp en kvast framför ett julgransträd.
Pojke i röd pyjamas med pingviner och snöflingor på dem spelar en Pokemon kortspel.
En man i kostym underhåller fyra barn.
En blondhårig kille i röd skjorta som rider.
Två kvinnor tittar på kameran leende sitter i stolar.
Ett blond huvudbarn som går med ett rött papper i handen.
En unge med en grön hink över huvudet.
En brunhårig kvinna håller en pojke i en skjorta med Reindeer på och en kockhatt.
Barn i rött under julen tittar på Toy Story leksaker.
En äldre dam sitter bredvid en bokhylla medan hon försöker underhålla ett litet barn.
Två små pojkar springer från en sjö med ankor
En Afrikansk amerika kvinnor i en hoppande hållning med hennes armar utspridda öppna och pyramidliknande strukturer bakom här
Barn som spelar fotboll på en plan.
Ett ungt gossebarn i gul skjorta som matas med en banan.
Två unga pojkar som lagar mat i ett kök.
Ett lyckligt barn med en Elmo-tröja i baksätet på en bil.
Tomten och mrs Klaus poserar med ett litet barn.
Ett litet barn besöker med någon klädd som en Disney karaktär.
Ett barn som bär en Elmo t-shirt står i tomtens släde.
En liten pojke sitter i en bil på en åktur.
Ett litet barn sätter en prydnad på en julgran.
En pojke blåser ut ett ljus på en tårta med en pingvin märkt "Grattis på födelsedagen, Quinn."
Ett litet barn i en röd overall står ovanpå en present.
Ett barn som bär en skjorta dekorerad med Elmos ansikte håller en röd ukulele.
Person mitt i ett ramphopp.
Ett spädbarn med mörkt hår som badas i ett litet handfat fyllt med tvålvatten.
En gatumusiker spelar trummor i en tunnel.
En grupp människor som sitter på stranden med en hink musslor.
En man som öppnar bakdörren till sitt parkerade fordon längs en sandväg.
Mannen som passerar dörren bär en vit skjorta och svarta löparbyxor med vita ränder på sidan.
En flicka i färgglada kläder på stranden
En snowboardåkare är silhuetterad mot solen när de lämnar marken.
Folk njuter av en måltid tillsammans under semestern.
Ett litet barn går längs en sjö med ett stort vitt tält i närheten.
Två småbarn sitter i en färgglad playpen.
En pojke som gör ett cykeltrick är i luften och väntar på att komma ner igen.
En brottare kastar en annan brottare till marken.
En man tar en tupplur på trottoaren i en upptagen stad.
En liten pojke i en röd jacka som utforskar en stenig terräng.
En person på en gul snowboard gör några tricks i snön.
Två små barn leker med leksaker.
Två unga flickor med huvuddukar står nära en dörr medan man läser en bok.
En skäggig man cyklar på stranden.
En man som är krökt på en klippa tittar på havets lugna vatten.
Lilla flicka som äter en suger mellan två bilar.
Folk i ett rum med blå färg och en dörr ovanför huvudet.
Pojke som gör en muskel håller papper som säger påskägg jakt.
Ett barn som leker med bubblor och går.
Två män seglade i en motoriserad flotte-typ båt.
En man håller upp en orange sjöstjärna medan han står i bröstet djupt i havet.
En man leder en grupp barn utanför hemmet.
En man med solglasögon och mössa håller i ett litet barn.
En kvinna med hatt som pekar ut i fjärran.
En basketspelare i luften som ska göra ett skott.
En jättestor reklamtavla av en mans magmuskler
En man sitter i förgrunden, och en kvinna med en drink är i bakgrunden.
En cykelförare hoppar från en ramp.
En motorcyklist som kör fort på en väg på en grön Kawasaki-motorcykel.
En asiatisk pojke skålar när han spelar bowling.
Två manliga brottare mitt i en match.
En man och en liten pojke sitter och vilar mot en stenmur.
Två kvinnor med huvudkläder som tittar på varandra i ett offentligt område.
Mannen står på hörnet och spelar musik.
Fyra barn bredvid ett blått hus går nerför en gata.
En grupp barn sitter på en vägg.
Ett par afrikanska barn bär ballonghattar och stirrar på något.
Någon surfar på en jättevåg.
En man bär en tallrik mat på en gatuförsäljare.
En brun hund för tillbaka en boj från havet.
Två kvinnor klädda med halsdukar över huvudet ser argt på fotografen.
En liten pojke i gula kläder som springer mot ett blått hus.
Tre människor är nära ett träd och kvinnan rör vid ett av männens ansikten.
En kvinna springer ut i en blå rock.
En fotograf sitter på sin kameraväska på stranden.
En asiatisk man kikar genom ett skyltfönster.
En tjej fotbollsmatch med ett lag i rosa, den andra i ljusblått.
En tjej som böjer sig bakåt och håller i hatten.
En liten pojke flyr från havets annalkande vågor.
En cykelcyklist hoppar backen på sin cykel.
Ett litet barn rider nerför en snöig kulle på en röd släde.
En hund med en boll i munnen som sitter utanför.
Tre män med matchande skjortor, byxor och hattar och en man i morgonrock är i ett rum.
En musiker som håller i en gitarrfilm spelar in lite action.
En flintskallig man i svart Enrolling Stones T-shirt läser en bok.
En man i svart skjorta sitter i en stol.
En vit man spelar gitarr i en inspelningsstudio.
Musik sätts ihop i en studio.
En man står framför en motorskoter och håller upp en bild.
En person som utför ett snowboard trick på ett högt berg.
En grupp kvinnor håller ihop för att fånga en boll.
Folk är ute på natten.
Den lilla pojken står mitt bland fåglar som har samlats på trottoaren.
Folk som står i en byggnad och tittar uppmärksamt.
En man som bär en Enrolling Stones t-shirt spelar på sitt Yamaha-tangentbord.
En skäggig man med ett tecken.
Två män sitter i kontorsstolar och tittar på en bild på en stor skärm framför dem.
En man klädd i grönt i en inspelningsstudio.
En stor grupp kyrkokörsångare på balkong.
Fyra människor skrattar och sitter på en soffa.
Ett gossebarn i vinterrock på en rund blå släde i snön.
En skuggig hund dammad av snö slickar näsan.
En person kastar ett föremål när en lurvig hund hoppar för att jaga det.
Tonåringar som maler en bänk på en skateboard
En man i svarta badbyxor dyker ner i vattnet
En man i uniform som delar något med en grupp barn.
En soldat och religiösa präster som undersöker och lägger ut bönemattor.
Två stora måsar är i vattnet.
Ett barn kommer ut ur ett rörglas och är på väg att träffa sanden.
En man och en kvinna som poserar framför ett julgransträd.
En grupp människor omger ett gäng uppblåsbara rosa stjärnor.
En boxare hoppar i snön.
Åtta medelålders par dansar och sex andra människor minglar på dansgolvet som ett tremannaband bestående av en gitarr, banjo och dragspel på en scen.
Den här mannen är klädd i vitt.
En man med skägg i grå skjorta som tittar i spegeln och rakar huvudet.
En man pratar på sin mobil i en stad.
Två män utför kampsporter, de är klädda i vitt och en man har sitt ben mellan benen på den andra mannen.
En man hukar sig på marken.
En man och en flicka som går på stranden, orange solnedgång bakom.
Två gamla män står nära ett bord i en McDonalds.
En brun hund med svart krage som skäller i snön.
Två fåglar interagerar i gräset
En stor vit hund är på väg genom ett snöigt fält.
Två män och en kvinna interagerar vid ett bord.
En man och två kvinnor har ett livligt samtal på en fest.
En kvinna som sitter vid ett bord framför tårtan.
En man och kvinna sätter födelsedagsljus på en tårta.
En fågel som plaskar runt i en bäck.
Fyra flickor hoppar upp och ner på sanden nära havet.
Man i brun skjorta på solig gata, en publik i bakgrunden
En kvinna med halsduk pratar med en man i glasögon.
Här är ett gäng människor som njuter av middag och chattar.
Tre leende människor och två andra inte vända kameran står utanför ett skjul på natten.
En grupp människor kommer att få sin fest på.
Tre små pojkar leker i ett stort snötäckt fält
Två män klädda som Santa Claus uppträder i en park.
En man håller ett pro Judéen protest tecken på en protest rally
Campare som sitter vid vattenbrynet.
Barn leker i gräs på en fullsatt utomhusfestival.
En man tittar över en liten klippa.
En blondhårig dam sitter vid ett skrivbord med en gul karta hängande på väggen.
En ung man som hoppar på ett rött räcke
Ett litet barn försöker balansera på en bänk i parken.
En kvinna går utomhus nära en kanal.
En grupp på fem män står mitt i ett rum som faller sönder och överges.
Ett kvinnligt patent på ett sjukhus som sticker ut tungan.
En pojke som bär en blå hjälm cyklar med fötterna på styret.
En stor, svart hund övar på att attackera en brottsling på en uniformerad man.
En hund är på väg att få en godbit i munnen.
Folk pratar och besöker på en buss.
Ett danspar som dansar på ett dansgolv med strobeljus som blinkar.
En dam som dansar tango i rött och avslutar sin rutin.
En liten pojke i rött står ovanpå en sten med ett leende och utsträckta armar.
Cheerleaders klädda i rött och svart håller två hejaklacksledare över huvudet.
En man i röd topp och hatt som spelar vad som verkar vara ett musikinstrument.
En pojke kastade käppen med eld.
Tre män jobbar med att bygga på natten på en gata.
Svarthårig mogen kvinna sitter bredvid ett bord av produkter.
Tre män klädda i centuriondräkter sitter framför byggnaden.
Ett litet barn med gröna goggles lutar på ett steg.
En blond pojke torkar näsan på sin ljusblå skjorta.
Folk klappar medan två kvinnor leker.
En man i blå skjorta som tar en tupplur.
Tre hundar springer i snön.
Den svarta och bruna hunden ligger ner med den mindre hunden hoppar över ryggen.
En grupp män som springer på ett fält.
Det är två personer som går i sanden.
En man med indianväst som spelar trummor.
En grupp leende tonåringar sitter vid ett bord medan de spelar ett brädspel.
En brun hund hoppar upp i luften.
Tre hundar springer runt i snön.
En brottningsmatch slutade precis och förloraren är upprörd.
En pojke som sitter på en dinosauriestol och håller ett blått föremål.
En man med en röd hjälm i bergen
En brun hund bär en käpp i munnen över en istäckt damm.
En man gör ett trick med ett svärd och släpper in svärdet i halsen.
En cyklist utför ett hopp över ett vitt räcke.
En liten flicka sitter på en bänk med armarna ihopvikta.
Två unga damer sitter på en liten vara i skumma klänningar.
Två män går längs en våt gränd.
I poolen omgiven av växter, en leende flicka med en hink stänker en annan flicka.
En familj som poserar vid manteln och julgranen.
En collegestudent diskuterar när han bär glasögon, som om han är vetenskapsman.
En kvinna som spelar akustisk gitarr med mikrofon
Ett litet barn med blont hår, bär en blå skjorta och jeans går i skogen.
Två personer på väg ner för vattenflödet, kajakpaddling.
En man som står vid en båt vid en brygga omgiven av stenig terräng och vatten och två andra båtar.
Två hundar i randiga tröjor slåss i snön.
En muskulös man i en Speedo och en kurvig blondin i bikini går tillsammans på stranden.
En person går i vattnet med ett nät.
Vattnet sprutar på barnet med ansiktet genom ett uthugget hål.
En flicka i lila skjorta har en kudde.
En man med motorsåg snider trä till en staty av en man.
En kvinna hoppar ett hinder på en bana.
En person står bredvid ett stenmonument med handen nära huvudet.
En man sitter på toppen av ett berg.
En snowboardåkare glider längs en ramp över en snöig lucka.
En man använder en stor stolpe för att ta bort bokstäver från en skylt.
En gyllene hund passerar en blå boll till en annan gyllene hund på stranden.
En förälder som hjälper sitt barn att gå i snön.
En kvinna ler mot den skäggige mannen som sitter i fåtöljen bredvid henne.
En blond kvinna och en flintskallig man som sitter tillsammans.
Kvinnan skrattar när hon blir slickad av en brun hund.
En person som dyker i en kelpskog.
En familj går uppför stentrappor i en park med grönska överallt.
En skara människor som står i träd.
En man håller i en mikrofon medan hon uppträder med sitt band.
En kille med en kvinnlig insektsdräkt på.
En kvinna gör ett handstånd på ett blankt golv medan två andra står i närheten.
En kvinna som bär huvudbonad och håller ett spädbarn
Två män, som är tvillingar, bär matchande svart skjorta och är på väg att slåss.
En kvinna går med sin stora väska.
En ung man visar sin spänning vid ett utomhusevenemang på natten.
Två vuxna och ett litet barn ställer sig utanför en bostad.
En äldre man sitter på ett tak och håller en hammare.
En man i grön skjorta håller på att fixa en cykelkedja
En vit kille med blå shorts på väg att slå en tennisboll med ett racket.
En man klädd som tomten sitter på en stol och spelar banjo.
Den här unge mannen bär en svart keps och klänning, och han håller på sin keps.
En kvinna rullar färska tortillas.
En man med hjälm gör ett stunt med sin BMX cykel.
Två kvinnor handlar glas utanför en butik.
En hund går i en däckbana i snön.
En kvinna går nerför en livlig gata och bär på papper.
En kvinna med en Nike hatt hårt på jobbet.
En man i jeans och en t-shirt som lastar något i en husvagn.
Afrikanska människor går förbi en tölfärgad byggnad i öknen.
En man cyklar längs en grusväg.
En afrikansk kvinna går bort från gräsiga hyddor i en by som bär en rygg i sin vänstra hand.
Människor från en afrikansk stam samlas utanför.
Deras ryggar mot kameran och under artificiell belysning står tre män vid matdisken.
En kvinna i vit och orange klänning dansar med en man.
En man står i ett gathörn och ett litet barn tittar på en skylt.
En militär grupp står i centrum.
Afrikanska människor i stamkläder i en öken.
En afrikan går genom ett fält.
Ett stampar poserar för en bild och mannen håller ett gevär på axeln.
En livlig stadsgata full av människor.
En närbild av en man och en kvinna.
En person bär en snowboard över djup snö.
En man som bär hängslen gör en split i luften.
Två bruna hundar leker i snön.
Mannen i den svarta jackan går förbi de förfallna dörröppningarna.
Flera människor spelar och koppla av på stranden.
En förare blir hög i luften med sin motorcykel.
2 kvinna bredvid ett bord säljer olika saker
En svart hund och liten vit och svart hund tittar upp på en köksbänk.
Fyra personer och en hundlek i snön.
En nygift hustru är under ett paraply som hålls av en pastor.
Män som bär förkläden arbetar i köket.
En försäljare tillagar mat finns det två röda gasburkar med mat på rad redo att sälja.
En man surfar på en enorm grön våg.
En dam med vänliga ögon och långt brunt hår håller en yxa vid ett träd.
En dam sätter fast någons skridskor i snön.
Fyra tjejer i blått uppträder på en basketplan framför en publik.
Cheerleaders, bär blå skjortor och svarta shorts, dansar i ett gym.
Två män brottas medan andra tittar
En man i blå rock med ett tecken.
En hund som ligger ner på en grön kudde.
En ung pojke håller i en tidning, som säger "Radeo", ovanför sin hemmagjorda radio.
En kvinna med långt brunt hår står utanför i snön och håller i en harpa.
Kvinnan med blont hår poserar med en stor yxa.
En kvinna håller två fans, en svart, en röd, och bär att göra med en röd klänning.
Två män i en grupp tittar ner på något.
En flicka sitter på en annons och kollar sin telefon; en annan flicka väntar.
Fem kvinnor som bär halsdukar på huvudet pratar.
En grupp människor är i en stor flotte på hackat vatten.
En stor skara människor som åker skridskor utomhus.
En kvinna leker med långa röda band på ett tomt torg.
Gamlingen tar en promenad längs de vackra böljande gröna kullarna.
En hund springer över en öken med buskar runt sig.
Den svarta hunden biter lekfullt den gula hunden nära möblerna.
Flera personer står och chattar i ett rum med många tomma stolar.
Många människor springer längs en gata i ett maratonlopp, som åskådare tittar på.
En liten flicka som sitter i en stol och håller en mobiltelefon i örat.
En person som bär orange rock går under mörka timmar.
En mans kraft tvättar trapporna vid en stor simbassäng.
Ett foto av en Volvo-återförsäljare på natten med två personer omgivna av apelsinkottar.
En pojke som bär röd skjorta stänks av vatten.
En äldre man som går på en gräs idrottsplats.
En person som bär jeans och en rock joggar på en trottoar.
De här människorna har trevligt.
En man ler när han sitter i ett bubbelbad och viftar med tårna framför kameran.
En stor man, i en jacka och hatt, håller upp något mot örat.
Musiker spelar nära en betongvägg.
Män i kostymer och slipsar som går nedför trappan
Flera personer klädda i rött sitter och står på gräs.
Ett passionerat, vackert, ungt par redo att dansa.
Fyra personer och en hund är på kanten av stranden.
En man tittar genom ett teleskop på något långt under honom.
En asiatisk kvinna som håller i en asiatisk baby som sträcker sig mot kameran.
Ett par tar ett bröllopsfoto med sin bröllopsfest.
En ung kvinna i en rutig jacka och ansiktsmask kör en passagerare på en skoter.
En skateboardåkare utför ett stunt.
En slalomåkare som bär röda byxor och svart skjorta åker förbi en röd flagga.
En skidåkare som åker nerför berget.
Två män på stranden med eld i ändarna.
En person som ritar kinesiska tecken med fötterna.
Tre unga flickor, som ser ut som systrar, håller alla rosa och blå baseballhandskar och en baseball.
En liten flicka som sitter i snön
Två killar poserar med två kvinnor, alla bär svart och vitt.
Vit, långhalsad fågel med gula ben flyger över vatten.
Unge man som flippar av något i en vattenförekomst.
Tre skolbarn i uniformer hopprep
En man i kamouflagejacka som drar en liten flicka i en ljus lila jacka med rosa mössa på en släde genom snön med en ATV.
Det finns en kvinna som bär en boll och ler.
Gymnast gör en volt över baren.
En brud som gör sig redo med sina tärnor klädda i rött.
Mannen rider en stor våg på en surfbräda.
Brudens sida av en bröllopsfest.
Två skidåkare gör sig redo att hoppa av en skidlift.
En man surfar över en enorm våg i havet.
Kvinnan i rött knäböjer för att hjälpa sittande bruden sätta på sig sin sko.
De unga vuxna står utanför skolan.
Två brandmän, klädda i uniformer, går ut ur brandbilen på trottoaren.
En person står i ett vidsträckt fält av smältande snö.
En skara människor står framför en stor byggnad med blekmedel framför sig.
En schäfer springer genom snön.
Pojke hoppar i luften med en skateboard.
En grupp synkroniserade simmare.
En man som romantiskt kysser en kvinna på en parkstig.
En man i Texas Longhorns hatt använder en spikpistol på taket.
En enda man i en blå t-shirt, jeans och en basebollmössa arbetar på ett tak i ett hus med bältros.
Ett barn i vit och ljuslila kläder som gråter.
En kvinna i en blå jacka får en cigarett utanför.
En rodeo-kille i röd skjorta rider på en bronco.
En takläggare i grå tröja och orange hatt går på ett ofärdigt tak vid ett sjönära hem.
En skogshuggare hugger ner en stor trädstam i karga skogar.
En folkmassa skriker utanför en byggnad som viftar med amerikanska flaggor.
Tre män sjunger med två mikrofoner.
En man i svart vinterjacka och röd skjorta står över en snöig sluttning med bergen som bakgrund.
Grupp av vuxna som sitter i en cirkel på ett möte.
En kvinna i en puffig röd jacka poserar för en bild på en skridskobana.
En grupp män, kvinnor och barn.
Surfaren kommer in från en stor våg.
En ensam snowboardåkare som hoppar i luften och gör ett trick.
En grupp på fyra personer går nerför en snöig gata.
En man ger ett barn till en annan man när de lämnar en båt
En liten vit och svart hund hoppar över en stor brun soffa.
Ett barn i vit skjorta och hatt klättrar.
Den svarta hunden hoppar ur snön för att fånga ett föremål.
En enda person ro en liten båt på en sjö.
En man dumpar en svart soptunna full med skräp i en maskin.
Vissa människor i byggnad som setts från gatan på natten.
En grupp människor som går på sidan av en järnvägsbana.
En man hoppar sin smutscykel på natten.
En urbefolkning som stod på stranden och skrattade åt fotografen som tog bilden.
En pojke sitter i en kundvagn.
En grupp klättrare i silhuett stirrar mot solen över bergstopparna.
En stor grupp människor står utanför en byggnad.
En liten hund bär en grön tröja och en ryggsäck går genom snö.
En man beundrar konst på ett museum.
En kvinna som bär en vit hatt som håller en lie och en skärning av vete.
En gentleman som häller upp ett glas vin till en dam.
Två män sitter på svarta läderstolar, och en av dem håller upp en koffeinfri Coca-Cola.
En man breakdances på huvudet mitt på dansgolvet.
En pojke i brunt springer på en grusväg.
Surfer är mitt i en enorm våg.
En äldre man med vita topphat dansar med sin fru på en sammankomst.
En brun och svart hund som hämtar en blå leksak.
En grupp asiatiska barn är en del av en publik som sitter på blå bänkar.
Tre tävlingshundar springer för att avsluta ett lopp.
En leende man som bär glasögon håller ett gråtande barn i ansiktet.
En traktor dekorerad som en flottör för en parad
Två svarta män poserar för en bild med vinterkläder på.
En ung pojke som spelar piano.
En grupp män som stod runt med en kvinna i Japan.
En basketspelare med boll och försvarare.
En kvinna håller en träram i pool av vatten, som är på en snöig plats, och det finns 2 fler halvnakna män bakom henne i poolen.
Ett ungt par gör yogapositioner framför en toriiport.
En kvinna i vit tröja går förbi affärer längs trottoaren.
En kvinna håller ett barn och ler för bilden.
Barn sitter framför en dator medan deras lärare instruerar dem.
Hantverksman arbetar med trä och en spikpistol.
En basketspelare dribblar bollen medan en annan blockerar honom och en tjänsteman tittar på.
Basketspelaren släpper basketbollen i nätet.
Det finns två kvinnor på hästryggen.
En man på en halv pipa som gör ett skateboardtrick.
Skateboardaren bär jeans och en vit skjorta utför ett trick.
En pojke och en person utanför kameran spelar ett kortspel.
En brun hund springer genom ett fält med öronen flygande i luften
En cykelförare i luften ovanför en ramp.
En äldre man som rakat skägget av en yngre man inför en folkmassa i en föreläsningssal.
Barn som bär svartvitt uppträder.
En grupp människor som sitter och står omkring på natten i kostymer.
Två barn hänger från en låg trädgren
En vit dam i färgglad klänning som dricker ur ett glas.
Två sumobrottare slåss i en match
Två sumobrottare slåss i en ring.
Ett litet barn med rött bälte gör en demonstration.
En pojke tar en tupplur när hans mamma bär honom på ryggen.
En man som sitter på en låda spelar gitarr.
En svart kvinna i vinterkläder som står i en byggnadsingång.
En man som korsar en korsning och andra går
Folk ser på när något lyser upp himlen.
En kvinna som rider på en barnleksak.
En trio av gitarrister, klädda i svart, spelar sina instrument.
Den här mannen gör ett stunt på en skateboard utomhus.
En man i grönt sparkar en fotboll medan en man i lila och vitt faller ner.
Det finns en massa människor på scenen som höjer händerna i luften.
En svart häst med vit på pannan och näsan, springande.
En grupp människor som hejar och roar sig.
En man i en blå nålstickad kostym läser en tidning medan han röker en cigarr
Kvinna i vit dribblande basketboll.
Sju barn sitter nära en person med svart blommiga kläder.
Unga män spelar fotboll på en strand.
Tre personer bär ögonbindlar med en Greenpeace skylt hängande i bakgrunden.
En dalmation går längs stranden.
Två unga pojkar som bär matchande New York Giants kläder leker med tvätt.
En ung person som leker i snön med två svarta hundar.
En grå terrier löper i ett snötäckt fält.
En skidhoppare är i luften.
En man med en namnskylt som säger "Jim" stickar.
En blond kvinna sitter under ett kalkongårdstak.
En skateboardåkare i luften högst upp på rampen.
En liten hund springer genom gräset.
Skateboardaren hoppar sin bräda i luften medan en annan skateboardare klockor.
En greyhoundhund sprintar.
Den vita och bruna hunden leker i det döda gräset.
Två män, en klädd i en blå nålstrippad skjorta, sjunger karaoke
En grupp kvinnor sitter runt ett bord och arbetar med garn i ett trångt rum.
En man som vrider en flammande batong.
Brun och vit hund leker med blå boll i blått vattenfyllda skal.
En kvinna och en man cyklar över en gata.
Det är många människor som trängs runt en blå skylt.
En man i orange håller upp en cykel nära en publik.
En liten vit och svart hund som jagar en något större brun hund i ett gräsbevuxen område.
Två personer i en orange racerbil.
Båten med passagerare lyfts upp ur vattnet med en stor kabel.
Barn som leker i vågor med solen vid horisonten.
En ung flicka leker på en skogsstock.
En mamma håller sitt barn på en röd soffa medan de båda har kul.
En man i röd jacka och hatt pratar med en annan man.
En pojke väntar utanför ett fönster med galler.
En skidåkare i röda byxor är på en snötäckt sluttning.
En grupp män dricker på en bar och pratar.
En kvinna sitter på ett heltäckningsmattat golv med ett barn.
Den bruna och vita hunden leker i snön.
En man, kvinna och barn sitter och äter mat utomhus.
Ett barn och en man som går i sanden.
Ett litet barn som bär en vit rock och spelar ett barnguldspel.
Tre personer poserar på sidan av ett berg.
En häger flyger genom luften nära lövverket.
En cyklist fotograferas när han hoppar från en ramp.
En man och en hustru står vid växeln när de gifter sig.
En man sopar gatan framför ett träd.
En kvinna som kysser en man i orange skjorta och brun jacka på kinden.
Två blonda kvinnor sitter i gräs med en liten hund.
En ung kvinna i gul skjorta löper över ett gräsfält i konkurrens.
En man står framför en krittavla som pekar på diagram
En hund tuggar på en metallstolpe.
En asiatisk man pratar på mobilen i sitt bås på jobbet.
Tre kvinnor springer med siffror på bröstet.
Flera personer pratar med läkare i ett rum.
En brun hund gräver lyckligt i sanden.
Två barn går uppför trottoaren med sina ryggsäckar.
Far och dotter leker i ett grunt område av en sjö tillsammans.
En stor fågel sveper ner mot marken.
Åtta män och kvinnor poseras med armar utsträckta i ett steg mode.
En grupp människor tävlar över ett gräsfält.
En pojke skateboard på en järnväg och tre pojkar tittar på.
En skara människor står på en snötäckt kulle och ser solen gå ner.
En vit och brun katt fladdermöss på en sliten sträng dinglande framför honom
En liten pojke som ligger på magen på gräset.
En grupp män i olika färger har ett maraton.
En ishockeyspelare tar vatten från en grön flaska.
En man med skidmask, klädd i svart, spelar gitarr.
En pojke i vita shorts står på ett rostigt torn.
En man förvränger sin kropp när han spelar baseball.
Man med muffins och kaffe överväger uttalandet "Vem är du?"
En man har somnat med munnen öppen.
En kvinna tittar på barn som simmar i en allmän pool.
Barn sover på mattor på golvet.
En hockeyspelare i blått och rött vaktar målet.
Två personer ler under en stor röd blomma och framför en vinvägg.
En man i grön rock som använder ett förstoringsglas för att läsa en bok medan han sitter på en bänk.
En kvinna som bär en vit jacka går förbi en skylt som annonserar hamburgare.
En man som bär en gul tröja bär en vit vagn på trottoaren medan en annan man som bär en ryggsäck går förbi.
En man är vid en shoppingvagn med folk som går på gatan.
En man med fyra löparhundar i naturen.
Ett team av breakdancers sätter upp längs sidan av en väg i staden när många åskådare samlas.
En fotbollsspelare i vit skjorta sparkade ett mål.
En man i vita byxor spelar gitarr, sjunger, medan två andra bandmedlemmar spelar med och dansar.
En man i grå skjorta sjunger på en mikrofon.
En man som spelar gitarr och signerar bredvid en kvinna i en klänning och spelar ett instrument
En man står bredvid en livräddare.
Tre personer spelar i ett band.
En kille med grå skjorta och jeans står på scen och sjunger med mikrofon.
En tonåring med en lila bandanna runt halsen spelar elgitarr och skriker in i en mikrofon.
Två unga kvinnliga innebandyspelare slåss om bollen.
En tonåring hugger ved på en snötäckt gata och en annan tonåring springer ut till honom.
Byggnadsarbetare som arbetar med virke med handskar.
En kille skär trä i små bitar i snön.
En snowboardåkare flyger genom luften.
Två personer cyklar på en ledig gata nära havet.
En kvinna som bär hinkar i bergen på landsbygden.
En leende man som lutar sig åt höger står bakom en leende kvinna som lutar sig åt vänster.
En man som rullade på en skatepark.
En surfare går upp en våg av vatten.
En man i en dragkedjad jacka snowboard.
En man i vit skjorta spelar tennis på ett fält.
En hund galopperar på stranden.
En man i hjälm står på motorhuven på en bil som brinner när folk ser på.
En far och en son som har roligt vid en pool.
En svart och vit hund bär en stor käpp på det gröna gräset.
En hund hoppar i luften för att fånga en frisbee.
En ung kvinna jobbar bakom disken på en juicebar.
En man som säljer kreativa ballonger på gatan.
En person som bär skidor hoppar över snön.
En person bowlar på en färgglad bowling allierad.
En man cyklar nerför en väg och följs tätt av en schäfer och möjligen en svart Labrador när två yngre män går längs trottoarkanten mot dem.
Två män talar nära på en fest.
En snowboardåkare som flyger genom luften och gör ett trick på ett snöigt berg.
Två kvinnor är i ett kök och lagar grönsaker i en wok.
Den unge mannen flyger genom luften på sin gröna snowboard.
Två människor (en man och en kvinna) lutar sig mot en byggnad samtalande
En kvinna som står i en grupp människor på ett kontor som en miljö.
Två gruvarbetare arbetar i en stor grop.
En svart och vit hund lämnar tillbaka en käpp i snön.
En man med vit hatt på en skoter.
En kvinna med rosa hår är ute med en grön rock och en halsduk med hjärtan på.
En snowboardåkare som får luft på natten.
En polis lutar sig mot sin motorcykel och tittar på gatorna.
Två personer på spjälsängar tittar på vattnet vid skymningen.
En person i röd skjorta på en skateboard.
Fyra asiatiska kvinnor poserar för en bild.
Folk har ett samtal i det inre rummet på ett skepp.
En person hoppar en cykel från en stor jordramp.
En grupp män och en flicka står på gatan.
Afrikansk kvinna med barn skriver alfabetet på en krittavla.
Två män för en diskussion på en trottoarkant medan en gul taxi kör förbi en kaotisk bakgrund av reklam.
Vuxna står runt ett klassrum i Afrika.
Folk samlas på en plattform i vatten för en ceremoni.
Barn spelar musik utanför.
En person gör en back flip medan andra människor och bilar går förbi i bakgrunden.
Ung rödhårig man spelar elgitarr.
Två vita hundar som springer på marken täckta med färgglada fallna blad.
En afrikansk kvinna klädd i traditionella kläder spelar trummor.
Byggarbetare använder en maskin på natten.
Dam i svart står och röker med en annan flicka som sitter på trappan.
Ett bergslejon hoppar från en klippa.
En skidåkare gör ett hopp med sina skidor korsade.
Två kvinnor stannar för att få sin bild tagen utanför chokladfabriken.
En dam på styltor på trottoaren har åskådare.
En äldre man sitter på en röd bänk med en yngre man.
En skallig örn står i grunt vatten.
En liten flicka i lila rock stirrar på fisken på marknaden.
En skateboardåkare utför ett trick på en ramp.
En blond hund fångar en boll i munnen i snön.
En familj på sex och tre hundar tar en promenad i skogen.
En grupp små barn som står i rad lutar sig mot en vägg.
Cyklist i snöig skog på natten
En kille är på marken i en tjurfäktning nära en halv luftburen vit tjur medan en annan kille går mot honom.
En person som står på styltor böjer sig över.
En vit hund med bruna öron springer genom snön
Ett litet barn leker på utrustningen i parken.
Två hundar springer genom en gräsbevuxen plats som är omgiven av träd.
En tjej får en tatuering på handen.
Två tjejer klädda med sumobyxor brottning medan folk tittar på.
En läderklädd rodeo cowboy stjärnor blankt, medan folk tittar på utanför ringen.
En grupp människor vandrar i skogen.
En äldre kvinna tillsätter kryddor till maten hon tillagar.
De matar sköldpaddsvattnet och pojken ser fram emot det.
En familj som bestämmer vad man ska göra på en restaurang
En snowboardåkare hoppar från en hög stenmur.
Två personer står bredvid en get.
Den nobbade hunden med nummer åtta lopp på grusspåret.
En kock använder en mikrofon när han öppnar locket på en ny maträtt.
En ung man med dreadlocks och en bunden färgad skjorta gör tricks på sin skateboard.
Nån i blå rock och vita sneakers är luftburna.
De unga vuxna tar en gruppbild av sig själva.
En person prydd i vitt kör en motorcykel.
Två små flickor, en i grönt och en i lila, läser en bok.
En pojke i blå skjorta springer medan han ler.
Man i blå och vit uniform skytte basket blockeras av man i vitt och rött.
Afrikansk amerikansk kvinna i blå skjorta tittar ner på mat.
Kvinnan med glasögon målar den blonda flickans ansikte.
En man ger gester till två kvinnor medan hon står på en parkeringsplats.
En vit man som bär vita och röda badbyxor hoppar in i en simbassäng.
Turister samlas framför en historisk byggnad på vintern.
En man i grå hatt skjuter någon typ av utrustning över isen.
En hund är bunden till vattnet.
Ett barn som bär grå vinterrock och blå snöstövlar är olyckligt när det upptäcker sitt lekhus täckt av snö.
Den här mannen studerar kontrollerna när han arbetar med tunga maskiner.
En man driver en liten utrustning.
En flicka med flingor i munnen.
En person joggar på en vattenkant i en röd jacka och svarta byxor.
En ung flicka rullar ut en jättestor snöboll.
En grupp människor går i dimman mot ett läskigt hus.
En flicka hoppar upp i luften framför havet.
En tjej i kostym dansar som andra tjejer i kostym.
Folk står och tittar på monitorer på väggen.
Folk syns knappt förutom upplyfta armar.
Många hundar visas i gräset.
En liten flicka blåser bubblor på en gård med ett skepp i bakgrunden.
En man kör en röd ATV uppför en oländig kulle.
En man med regnbågshår och en kvinna skriker ut genom fönstret på en limousin.
Många klättrar på en repbana utanför.
Mannen i ljusgul jacka och svarta byxor rider en cykel i snö på en väg som skyddas av ett räcke.
Killar i blå skjortor jobbar på en bil.
En ung man jonglerar sex svarta och vita bollar.
En medelålders kvinna, bär förkläde, bär en behållare med glass och kottar.
Mannen sitter på en pall och spelar trombon.
Tre hundar springer på bred, gräsbevuxen, utomhus område.
En hund i en sele som drar en rosa bärare bakom den på snö.
Ballerinas dansar på en stor scen under blå spotlights.
En man ligger mitt i en smutsig gränd.
Ett barn tittar på en snowboard i snön.
Skidåkaren lutar sig framåt i snön.
En snowboardåkare hoppar över en snöig kulle
En brun och vit hund står på sanden för att titta på en annan hund.
En performancegrupp iscensätts i en gemensam rörelse.
Stor svart hund drar runt saker på en röd släde.
Grupp av människor samlades för en begravning på en strand.
En man ristar ett isblock med motorsåg.
En äldre man som bär en klargrön, gul och röd skjorta som håller ett rött dragspel.
Cyklister tävlar i ett lopp som tar dem på en grusväg.
En hundsläde med två passagerare som färdas genom snön.
En brun ekorre hoppar upp i luften i ett snöigt område.
Tre fönsterbrickor utför sitt jobb.
En ung flicka med mörkt hår och en röd rosett ler samtidigt omfamna en ung mörkhårig pojke.
Folk står på en isig gata i snön runt en bil.
En deltagare i ett hundspannlopp passerar åskådare.
En liten pojke beundrar en grön sportbil.
En grupp människor är på ett konvent och viftar med amerikanska flaggor.
Tre hundar springer i jorden.
En man försöker ett trick skott i en liten bowlinghall medan hans vän tittar.
Killarna skjuter.
En liten flicka i randig klänning har en rosa halsduk.
Folk leker på en snötäckt gata.
En clown i svarta och vita randiga skjortor underhåller en ung flicka.
En äldre kvinna som sitter vid ett bord i en restaurang och håller i ett glas.
Två män jobbar på trottoarkanten.
Man ritar en bild på en balkong med utsikt över en kyrka.
En schäferhund springer i snön.
En pojke kör genom ett stort hjul.
Två pojkar springer i en metalltunna.
Två kvinnor med svarta väskor tittar på baksidan av en kamera
En man i tung rock reparerar på en tågstation.
Två vita vanliga pudlar som spelar dragkamp i snön.
En brun hund som håller en stor käpp i munnen och springer i snön.
En blå karaktär sitter i läktarna på ett sportevenemang.
En volleybollspelare i en orange skjorta hoppar upp i luften för att träffa bollen.
Två kvinnor i orange hoppa upp för att blockera en volleyboll skott på en volleyboll match.
Två bruna hundar som bär mynningar tävlar genom ett gräsfält.
Den leende kvinnan står i gräs nära en bäck.
En flintskallig man med brun jacka står framför Bryant Parks tidningsställ medan snöfloder faller på New York.
En grupp människor tävlar.
Folk framför en beige femvåningsbyggnad.
En man ligger på en säng och öppnar ett paket.
En kvinna i päls och hatt tittar på blommor
En liten flicka går längs den trädkantade vägen.
Tre personer är klädda i jadegrönt och pratar nära ett staket.
Folk tittar på konsten i utställningen.
Två snowboardåkare i gult och grönt hoppar i luften.
En man i en skogsmiljö tittar genom en ihålig träbit.
Två killar med långt hår som står framför ett fönster.
Ett pojkbarn håller i en fladdermus som han ska svinga mot en pinata.
Två unga män står vid ett hems öppna ytterdörr en snöig kväll.
En grupp på fem vuxna ställer sig framför byggnader.
En mamma är på knä och lagar sin dotters blå klänning.
Mor och dotter åker upp till stan för att shoppa
En skidåkare som bär vita solglasögon åker nerför ett snöigt berg väldigt snabbt.
Medelålders man som städar den fallna snön på taket på sin bil med en kvast.
En flicka i svart rock och röd hatt rider en röd släde nerför en snöig kulle.
Två unga barn som bär vinterrockar leker i snön.
En liten pojke berättar en hemlighet för en liten flicka
En sångare sjunger in i en mikrofon.
En brun och vit hund som går i snön nära ett staket.
En man går genom eld.
En man på marken nära en rad bilar, och en annan man som står och håller den första mannens ben.
En man som hoppar från några stockar.
En kvinna kollar hur det går med avläsningen av ett löpband på gymmet.
En man i blå skjorta vandrar genom en naturstig.
En person sitter på en strand med regnbåge i bakgrunden.
En grupp damer som spelar kort
En kvinna knuffar en barnvagn förbi ett staket bakom vilket några uniformerade pojkar sträcker ut sig.
Två män tävlar i vattnet.
Flera surfare är ute i havet och väntar på en våg.
En pojke och en ung kvinna i en huvudduk gör fredstecken.
En svart och vit hund som hoppar i snön.
En ung flicka leker med sina dockor.
En brunhårig man med glasögon bär en bourgognetröja medan han sitter vid ett middagsbord och kollar sin mobil.
En man och en kvinna sätter upp en kamera.
En liten flicka i en rosa jacka är i mitten av ramen.
En man intervjuar en pojke i en samling människor.
En man är uppslukad av lågor medan två filmbesättningar övervakar.
En man som spelar gitarr och en man som spelar trummor
Grå hund med mynning och med # 8 gul randig identifiering körs.
En kvinna med mörkt hår som arbetar med färgstarka tyger.
En svart hund med lila krage och ett svart koppel springer i gräset.
Vackert bergslandskap och skidlift.
En grupp ligger i snön medan någon på en blå snösläde hoppar över dem.
En man som dansar på gatan inför en folkmassa.
En man sätter upp en kamera på ett stativ medan en kvinna står i bakgrunden.
En man som sitter framför en scen
En kvinna i svart rock med en kamera på ett stativ
En man spelar gitarr framför en tegelvägg.
Ung pojke i en vintermössa som glider nerför en snöig kulle.
Mannen i vitt spelar basket mot mannen i blått.
En solbränd och vit hund går i sanden en fin dag.
En hund springer rakt mot ett hinder.
En hund tittar på en vit svan som simmar i en sjö.
En man står på huvudet framför en folkmassa.
En man som poserar framför folk på en livlig gata.
Man i färgglada jersey och mössa utför för publik i urbana området.
En pojke som springer genom surfing på en strand.
Två hundar springer över gräsfältet.
En man i svart skinnjacka somnar på kollektivtrafiken.
Flera barn springer tillsammans med en kvinna.
Folk samlas under färgat ljus i ett stort tält.
En man i orange snödräkt är på en hundspann i snön.
Hundar drar en person på en släde i snön.
Man i vit skjorta står framför vitt staket och stor byggnad.
En rödhårig flicka ligger i badet med suds över hela hakan.
Killen i svart uniform dribblar basket bort från killen i vit uniform
En gul plyschleksaksdräkt på gatuevenemanget.
En grupp män leker rugby.
En gammal vit man som spelar saxofon när han sitter på en pall.
En man koncentrerar sig på sin musik och håller i sin fiol.
Arbetaren står på en stege på en trottoar i staden och reparerar byggnaden med en stor borr.
Två fäktare i växelslagsmål i en fäktningsklass
De två männen spelar Frisbee på ett fält.
Två män lösgör sina nät på bryggan.
De två unga pojkarna leker i en pöl en skön dag.
En man håller i ett barn som håller i glasögon.
En person på en cykel hoppar högt i luften på en strand.
Flera barn sitter ner och håller basketbollar
En kvinna med en vagn med ägg går på en marknad.
Räddningspersonal hjälper en person in i en bärbar apparat, i ett snöigt område.
Unga asiatiska elever ler och presenterar sina nya basketbollar.
Ung flicka i rosa skjorta med leksaker runt omkring henne.
En räddningsman leder en man som drar en släde med nödutrustning på en snöig stig.
En svart och vit hund som biter på en bit is.
Tre personer står på scenen och två av folket tittar på när den andre spelar trumpet.
En ung pojke leker i parken med sin mor.
Två vita hundar simmar ansikte mot ansikte i skuggigt vatten.
En man med strålkastare står i en grotta.
En motocross cykel rids längs en skogsstig.
Två löpare gör sig redo att tävla på ett spår.
En gul hund springer nerför en grusväg.
En grupp musiker på scenen som spelar musik.
En motor-cross ryttare i rött stänker genom lera och regn med sin motorcykel.
En kvinna verkar kämpa för att lyfta ett föremål.
En vit hund med en orange fläck hoppar genom torkat gräs.
En pojke slipar en avsats på sin skateboard.
Folk i en pool och något skapade bara ett stort stänk.
Den bruna och svarta hunden springer över snön.
En mans himmel på den snöiga marken bland träd.
En man, i en blå skjorta, lyfter en vikterob.
En grupp människor skjuter upp en varmluftsballong.
Tre hundar tävlar i snön tillsammans.
En hund springer längs med en ko på ett gräsfält.
En hund och en kyckling bredvid en byggnad.
En kvinna i jeans och en svart jacka som står på vägen framför en vit och röd buss.
En man styr en blå båt förbi färgglada hus.
En brun hund som gör ett roligt ansikte medan han står på stranden.
En pojke på en snowboard hoppar genom luften.
En stor grupp människor packas tätt in i ett tåg.
Två personer är sumobrottning.
Lite svart hund och en stor brun hund är ute i snön.
En man som pratar med två kvinnor.
En svart kvinna och två svarta barn sitter i ett halmtäckt tält.
En parkeringsplats fylld med cyklar och trikes.
Ett kylskåp sitter fast i snön, och en man åker skidor på den.
Grupp av svarta män som lastar bagage på toppen av en buss
En kvinna i en lavendel tank topp säljer vattenkokare korn i en monter.
Flera människor sitter på ett tak i en stad i Mellanöstern.
Mannen sjöng en sång medan en annan man spelade gitarr.
Män som jobbar på ett projekt.
En man med orange skjorta träffar en boll med tennisracket.
En lättklädd man som har ett samtal med en man i kostym.
En man som är på väg att slå en tennisboll med ett racket.
En äldre gentleman sitter bakom en kontrollbräda.
En städerska i vit uniform sopar golvet.
Motocross ryttare hoppar sin smuts cykel.
Två flickor stod inne i en trägrind med en tjej som vinkade.
En violinist och en sångare uppträder inför folk.
En man som står och tittar på en bok och en pojke sitter och håller i något.
Man i blå skjorta rökning
Mannen spelar akustisk gitarr medan de andra männen gör gester
En motorcyklist som rider övertäckt huvud mot tå med lera
Tre kvinnor och män säljer sina varor på en kall vinterdag.
En grupp män som drar rep på en klippa.
En simmare kommer upp över vattenytan för att få luft.
En man sitter vid en dator och typer.
En äldre vit man med en blå hink som målar en fönsterbur.
Tjejen i skolan klär sig på toppen av ett träd.
En man dyker ner i vattnet nära en strand.
En mängd olika människor på baksidan av en stor vagn.
Två stora hundar springer medan en tredje klockor.
Tre kvinnor ler med målningar bakom sig.
En hund nipper vid benet på en häst.
Fyra unga kvinnor som bär bikini spelar beach volleyboll
En kvinna i formell ridutrustning rider sin häst på stranden.
Olika personer såg genom ett tunnelbanefönster.
En man i en bast och tunn mustasch gester till två kvinnor i samtal.
En kille på en skateboard som ska göra ett trick
En man som gör breakdancing på huvudet med en silverhjälm och en annan spelar musik medan åskådare passerar
Mannen bär flashig guldskjorta stående i lägenheten
En basketspelare försöker sikta på målet samtidigt blockeras av andra spelare.
Man gör ett trick som vänder över flera människor radas upp på en gata mässa.
En jordekorre står på kanten av ett fält och en väg
Ett par vandrare korsar en bro.
En liten brun hund springer i snön.
En smutscykel sliter upp terrängen.
En ensam skidåkare går nerför en tom kulle under en blå himmel.
Vit far och sol i blå våtdräkter med boogiebräda i vattnet.
Folk står på en järnvägsplattform och läser tidningar.
Folk i ett gymnasium dansar i en tävling.
Racinghunden har en munkorg och bär randig tröja #8.
Gubben har en röd skjorta på en grön bänk.
Tre män står tillsammans med två par skalor bredvid stora högar av färska grönsaker.
En vit kran flyger över lite vatten.
Två hundar springer genom gräs nära en vattensamling.
En rödhårig kvinna bär ett barn på bröstet i en bärare.
En man arbetar på ett mikroskop medan åtminstone fyra andra observerar och en videofilmar det.
Ett band som spelar i ett mörkt inomhusområde.
En man som bär halsduk runt huvudet spelar flöjt utanför.
En person som sitter fast i en sele svänger mot en upphängd boll.
Två hundar ligger på rygg på den lila sängen.
En man i röd skjorta håller i tidningar.
En man håller en hög med tidningar i en lobby, och en kvinna bredvid honom har tagit en av tidningarna och ler.
En ung flicka fyller en flaska med vätska med hjälp av en tratt och en kanna.
Ett barn i scoutuniform lägger saker i en affär.
Två män på ett kontor brottas när två andra vaktar.
Två personer som arbetar i vatten bredvid fält
Fyra damer i baddräkter spelar sandvolleyboll på stranden.
En man är uppe på en ställning och verkar tvätta fönstren i en byggnad.
En man med dreadlocks pratar på sin mobil.
En bebis i en blå skjorta som tittade på kameran medan de höll i en krita de använde.
En man och en kvinna som sitter vid vattnet.
En kvinna som täcker sina ögon i en park när dagen når sitt slut
En person i vinterkläder täcker sitt ansikte med en tröja.
Den bruna huvudpojken på sin skoter ska till leksaksaffären efter skolan.
En svart hund jagar en annan svart hund som bär en boll i munnen.
En krigskonstnär som visar sin skicklighet genom att bryta brädor med foten i en dojo.
Ett litet barn försöker hitta sin väg.
En grupp människor, varav flera bär luddiga rosa antenner.
Flera personer hjälper till att flytta en försäljare vagn.
En svart hund och en brun och vit hund som springer i gräset.
En grupp människor viftar med små amerikanska flaggor med ett staket.
Ingen trafik eftersom det är söndag och mannen väntar på att korsa vägen.
En svarthårig kvinna handlar mat med rosor.
Man i blå hatt och blå och svart randig skjorta gör skateboard trick på rock.
En man med rock och halsduk står nära ett café.
Ett barn med en pinne och ingen tröja sitter i gräset
Tre pojkar letar efter sina böcker i ett bibliotek.
Svart och vit hund hoppar upp i luften för att fånga en boll utanför.
Tre barn klättrar upp i ett stort träd i staden.
En hök sitter i ett spirande träd och tittar åt vänster.
Folk lyssnar på två män som spelar gitarr på en båt.
Flera människor går längs en smal bro över lite vatten.
Två personer vandrar uppför en snöig kulle.
En liten svart hund springer genom den vita snön.
Liten asiatisk man i shorts med en riktigt stor såghuggning trä.
Köksarbetaren på en restaurang observerar matsalen, inklusive en man i en röd jacka.
I en liten by sätter en man segel längs Swamp.
En frisör applicerar permed på en klients hår i en salong.
Två kvinnor poserar för en bild i ett sovrum.
En kvinna i en grå topp har sin spegelbild fångad i badrumsspegeln.
Två kvinnor och ett barn firar på en kvällsfest.
En individ går nerför ett steg med en väska i sin vänstra hand.
Två kvinnor brottas vid stranden bredvid en stad.
En halway har en skylt som säger "PORT DU CASQUE OBLIGATOIRE" och lite graffiti.
Kvinnor vid en disk i en tvättmatta tittar på genom hennes handväska.
En tonårspojke ger en annan tonårspojke en ridtur i skogen.
Valpar, kycklingar och en kalkon som undersöker innehållet i hinken på smuts.
Två hundar står och en hund ligger på rygg.
En affärsman åker tidigt för dagen.
En skäggig man i en blå skjorta skrattar medan en lämplig mustached man håller upp ett glas.
En man som tittar på landskapet genom kikare.
En man som är fäst vid en sele klättrar uppför en stenvägg.
En ung pojke utanför poolen, ler.
Den vita svanen lyfter från vattnet.
Två män springer med siffror fastsatta på sina skjortor.
Ett litet barn som bär jeans och en fotbollströja bär en klädeskorg som hatt.
En man bär ett nummer på sin vita skjorta.
Den här mannen verkar sova medan han vilar huvudet på handen.
En man som bär en maroonskjorta bunden runt ansiktet ligger på cementen.
Människan står framför ett bord fyllt med ett sortiment av ätbara föremål som mörker ser på.
Två afrikanska män sköter sig själva.
Sverals unga pojkar klättrar upp ur vattnet på en betong trottoar
En kvinna ligger på golvet bredvid ett barn.
En siluettfigur står på toppen av en snötäckt topp i slutet av vissa spår.
En man och en kvinna sitter vid ett bord med en drink.
Ett barn i rosa har ett föremål som verkar brinna.
En skateboardåkare hoppar från ett träbord nerför några trappsteg.
En cyklist som går uppför en stig kantad av byråkrati.
Ett barn sitter på en blå rutschkana.
En brun hund jagar en svartvit fotboll.
Gammal man och kvinna i jackor vända mot varandra
En lång snowboardåkare som hoppar över en barrikad utanför i snön.
Två basketspelare spelar i ett spel.
Två män spelar basket och en försöker blockera de andra skotten.
En basketspelare gör sig redo att skjuta en båge
En man på en sportslig även klädd i grönt och gult ler.
En person i en mångfärgad jacka som röker en cigarett inne på uppfarten till en byggnad.
En äldre vit man i svart cowboyhatt sjunger in i en mikrofon.
En svart hund springer nerför en stig.
Basketspelaren i blått löper mellan två spelare i vitt.
Basketspelaren håller bollen.
Den bruna och svarta hunden har sin mun öppen.
En hund i ett fält som håller något i munnen.
En kvinna i blommig skjorta och vita handskar balanserar en fiskbowl på huvudet.
Det finns hundratals människor med röda skjortor som springer ett maraton.
Två personer med skyltar som läser "Free Hug" stirrar med människor i närheten.
Folk som går nerför gatan kantade med kinesiska lyktor.
En man i grönt som håller ett tecken kramar en blond kvinna.
En kvinna med rött hår håller på med papper.
En kvinna och två unga flickor skyddar sig mot regnet med paraplyer.
Snöspolaren rider på en rail.
En kvinna gör yoga och ler mot kameran.
Man i en kontorsmiljö hoppar rep i affärskläder.
Två personer står framför en sjö i snön och poserar för en bild.
Två par poserar för en bild på vintern.
En stor grå fågel börjar landa i vattnet.
En flicka i Burka lär sig ordförråd i ett klassrum.
En tjej håller plastfolie runt huvudet.
En snowboardåkare går nerför en kort kulle bredvid trapporna.
En man med en röd vit och svart randig skjorta drar en vagn full av blå hinkar och kvast.
Några tittar på ett kryssningsfartyg.
En kvinna cyklar och njuter av havslandskapet.
En unge som sitter på en båt vid vattnet.
En flicka tröstar ett litet barn som föll på isen när hon åkte skridskor
En svart man med dreadlocks klappar.
Två svarta hundar springer med en tennisboll över den snöiga jorden.
En man i vit hatt städar ett skyltfönster på en restaurang.
En man som håller ett barn som klappar en ponny.
Två basketspelare som slåss om kontrollen över en boll.
En man i jeans och en arbetsskjorta och handskar håller en motorsåg med en växt i förgrunden.
Cricket spelare med röd mössa träffar bollen utomhus.
En man och en skateboard ovanpå en tunna.
Flera kvinnor spelar en omgång beachvolleyboll.
En pojke lutar sig mot ett baseballträ och håller ut en arm som är oåtkomlig.
Tre män bär blå hattar och orange västar.
En man som bär skyddskläder blir biten på armen av en hund.
Tre vänner skrattar på en skidresa.
Den lilla, gyllene hunden försöker ta ett lurvigt föremål från ett större utseende
En man med shorts springer längs en strand.
Inspektörer försökte kolla en bil som hade kolliderat med ett spår utanför Chevrons bensinstation i Texas.
En kvinnlig rugbyspelare som försöker outmaneuver motsatta spelare.
På gatan sitter en man och spelar trummor medan en man som står bredvid honom spelar gitarr.
Hunden springer i den djupa snön.
Unga flickor med guld och röda kåpor som springer i ett gymnasium.
Två personer är ute och går genom snön.
En man som bär en blå våtdräkt vaknar upp genom en stor våg.
Ett par delar en kyss en kall solig dag.
En moderiktigt klädd kvinna som håller en skiva i en ram i en begagnad bokhandel.
Folk samlas flygande drakar på en bergssluttning.
Den här personen ligger på golvet längst ner i trappan och saknar en sko.
En man som joggar på trottoaren när han lyssnar på musik.
En man skateboardar inför en grupp människor.
En man som gör en akrobatisk rörelse på havsstranden.
Hunden springer full fart genom ängen.
Servitris i svart hatt ställer upp bordet.
En man i våtdräkt surfar på en våg.
Person skidåkning på sluttning nära skidlift
Vita tält radade med röda kinesiska lyktor hängande från dem
Två hundar leker runt i smutsen.
Hunden står med 1 fot upp i ett stort fält.
En man på en bmx cykel hoppar över ett tåg
Ett stort fordon färdas genom en guppig och lerig stig.
En svart man går förbi en byggnad på en livlig trottoar.
Pojken är på blå cykel och är ovanför ett staket.
En man som går bakom en löparhund på stranden.
En vacker vit hund som går i det bruna gräset.
En grupp på fyra killar som bär tutu
En snowboardåkare spyr upp snö när han rider på brädan.
En bonde och tre barn arbetar på en gård.
En svart och vit hund vilar huvudet på en kamera.
En person med grön skjorta hoppar högt över gräset.
En liten brun hund leker med en boll på stranden.
Två flickor hänger tinsel från en julgran.
En tjej i svart skjorta sätter en stjärna på en julgran.
Två unga flickor är inlindade i julton.
Liten pojke med blå ögon bär en vit och röd, orange och gul haklapp
En liten pojke som skyfflar snö på uppfarten.
En kvinna går sin hund längs en rad färgglada hus med garage.
En man i vit hatt som tittar på måsar med två barn.
En kvinna i en svart och vit långärmad blommig printklänning med rosa läppstift verkar sjunga nära en tegelvägg och en atmmaskin.
Ung pojke i röd huvtröja skridskor.
En skidåkare hoppar från en brant bergssluttning täckt av snö.
En mountainbike som bär en färgstark hjälm rider nedförsbacke.
En man i alla svarta kläder på scenen läser något från ett papper till mikrofonen till publiken.
En del människor i medeltida kostym går genom en fullsatt gata.
Barn, småbarn och kvinnor som tar ett bad och tvättar kläder, förmodligen nära en flodbädd och en flicka bär en behållare med vatten.
En grupp människor står upp.
Tre färgglada clowner med ballonger poserar bredvid en annan plast clown.
Ett litet barn leker med hula-hoops på en gård i ett område.
Tre pojkar korsar en flod med något slags vilt djur.
En man med svarta handskar sitter på någons axlar för att ta en bild.
Tre män med vita uniformer står på ett gräsfält framför en folkmassa.
Asiatisk mor och barn tittar på akvarietanken.
En svart fågel i luften med löv i munnen.
Hockeyspelare med en chansning.
En kvinna i rött och vitt står mitt på gatan.
Pojke skateboard ner för en trappa räcke på vintern
En skidåkare klädd i svart hastigheter nerför berget.
En person som bär rosa byxor och en vit jacka är snowboard.
Tillbaka till en rödhårig kvinna som rider på tunnelbanan.
En pojke i blå jacka på ett tunnelbanetåg.
En grupp människor är på en båt i en marina.
En svart och brun hund springer med en tennisboll i munnen.
En kock i en blå hatt böjer sig fram inför folk medan de äter.
En ung pojke med ett blått paraply väntar utanför en affär.
Två kvinnor omfamnar, en i brun skjorta och en i lila skjorta, som andra människor ser på.
Barn som pratar med en äldre kvinna framför en dörr.
Tre barn står på en trädstam som har fallit.
Den här Gentleman i en vit skjorta, studerar verkligen, på sin dator.
En man sparkar fotbollen mot målvakten en varm dag.
En skidåkare klädd i rött på ett snötäckt berg.
En man som går nerför kullen i snön
En pojke med en basketboll.
En person i en grön skjorta på en skateboard hoppar från en kort uppsättning trappor.
En snowboardåkare i rött rider nerför sluttningen.
En kvinna i en överdådig orange klänning dansar med en man i alla svarta kläder.
Mannen leker på gården med två hundar.
Människor på cyklar rider genom en grupp åskådare.
Ett par njuter av ett glas vitt vin.
Tre basketspelare i vitt försvarar sig mot den anfallande spelaren med bollen i orange.
Fyra personer och solen.
En liten flicka som sparkar en fotboll till en liten pojke.
Ett barn gör några övningar för fotboll.
En grupp ungar springer medan de spelar fotboll.
En surfare i röd skjorta är under en stor våg.
En skakig svart och vit hund springer på gräset.
En man och en kvinna rider skoter som fordon
Ett barn som korsar ett kedjestängsel för att komma till vattnet.
En publikscen framför moskén.
En man som står ensam med en sorglig blick på sitt ansikte.
En man i randig hatt går förbi en discoanläggning.
Den färgstarka ryttaren rider nerför en kulle på en skoter.
En grupp cykelförare rider på gatan.
En kör står framför en amerikansk flagga i sjöman hattar sjungande.
En liten flicka i lila hatt står i huvudrollen.
Fem personer i vita skjortor med grå hattar i skogen med verktyg.
En pojke springer på färgstarka linjer.
En kvinna sover på en stol på en buss.
En tonåring försöker sig på ett skateboardtrick i ett stadsområde.
En liten pojke med blå glasögon och headset bär en svart skjorta med ett nummer på och en grå shorts.
Ett barn i en gryta på en spis.
Ett barn som bär kappa bland några träd och roliga mönster.
En kvinna med en stickad mössa på ler nära en Domino Pizza skylt.
Ett barn i en brun, mönstrad jacka ligger på en soffa med en blå filt
En snowboardåkare hoppar högt över den snöiga kullen.
Fyra personer går längs sidan av en tegelbyggnad.
En mountainbike som bär vita lopp genom en sväng.
En leende kvinna och man sitter framför en mikrofon i en musikstudio.
En åkare utför ett stunt från en cementvägg täckt av graffiti.
Massor av människor på en trappa i en gammal tjusig byggnad för ett evenemang.
En grupp människor som går på snöiga steg.
En stuntman gör en cykel trick upp i luften medan fyrverkerier går runt honom
En brun gud slappnar av på en trottoar.
En stor grupp människor samlas för att tillkännage sin sak inför kamerorna.
Människor klädda för svalt väder, ivrigt väntar i kö.
Två barn ligger på en säng medan de leker med leksaker.
Asiatisk pojke sätter sitt huvud i en stor bubbla.
Folk samlas runt ett bord med mat och utanför en taxi wisks förbi.
En tonåring tar en risk genom att dyka på sin sida.
Två pojkar leker i vattnet nära en gammal byggnad och en båt.
Två latinos spelar instrument; en på violinen och den andra på harpa.
Hane bär brun skjorta som håller en mikrofon med ett uttryck för sång.
En grupp artister sjunger och spelar under strålkastarljuset.
Två personer sitter på en brygga bredvid varandra och tittar på solnedgången.
En man som sitter i hörnet och pratar på sin mobil.
En grupp av många människor som verkar sälja eller äta mat under ett tält.
En kille som spelar gitarr med "Vad som än krävs" skrivet på den.
Flera människor har satt upp tillfälliga läger bredvid en stor marmor stödpelare.
En scen uppförs på en stadsgata medan förbipasserande vakter.
En snowboardåkare utför ett stunt framför en skara åskådare.
Turister som tar en bild framför en byggnad.
Ett lag av fotbollsspelare i vita remsor löper runt kottar på en idrottsplan.
Tre damer står i ett rum som ser ut som ett arbetsrum.
En äldre man med en rutig skjorta tittar genom ett mikroskop.
Åskådare tittar som en snowboardåkare gör ett trick.
En svart ung man i en blå skjorta för en livlig diskussion med andra ungdomar runt ett bord.
En ung pojke som rör sig mot en gul boll.
Två kvinnor i hattar står framför åskådare, den ena spelar fiol och den andra spelar dragspel.
Ett klassrum fullt av män, med läraren på framsidan.
En man som bär en t-shirt som har "gnu" tryckt på den ger en teknisk presentation.
En pojke surfar på en våg.
Står och sitter jämnt med en rad av träd, två kvinnliga figurer vänder sig mot riktningen av en vattenkropp.
En tyngre man med blå skjorta och svarta byxor går nerför trottoaren i ett köpcentrum.
En tjur tar sig ut genom grindarna på en rodeo.
Människor i en båt som svävar ovanför vågorna.
En vit häger flyger upp i skyn.
En liten flicka springer över gräset mot träden.
En brun hund går i snön mellan några tallar.
Läraren hjälper sin elev att slutföra en del arbete.
Kvinna med glasögon, håller en kamera, nyanserar hennes ögon med händerna medan hon står i förgrunden av en havsutsikt.
En tonåring klättrar upp för en stenmur.
Två män som bär brottningsutrustning med huvudet pressat ihop.
Tre barn leker i det grunda havet.
Innan ett par beställer sin mat på en restaurang bestämmer de sig för att clowna runt för det andra paret som sitter med dem.
Biker hoppar från en ramp i skogen.
En man spelar ett stränginstrument som en del av en orkester.
En kvinna i konisk hatt arbetar vid en smal vävstol.
En man i brun jacka som går ensam uppför en trappa.
En färgstark lastbil lastar av i en sjö mittemot ett tältläger.
Stoppa actionram för en racer i en cykel race.
Tre pojkar med blå skjortor som ler för kamerafoto.
Äldre svarthårig kvinna som lutar sig mot kanten av en tegelvägg med hängande tvätt bakom sig.
En fotbollsspelare hoppar i luften under en match.
En familj på nio sitter fullsatt på en vit soffa och ler.
En svart pudel med en repleksak i munnen.
En stor grupp människor som deltar i ett evenemang med leverantörer och mat.
En svart hund hoppar genom snön nära ett stängsel.
En ung man övar på sitt elektriska Yamaha-tangentbord.
Tre barn leker med metallmöbler.
En afrikansk amerikansk kvinna cyklar nerför gatan.
Leverantörer säljer frukt och grönsaker på en utomhusmarknad.
En man går förbi en butik som har ett namn på franska.
Två unga vuxna ler mot kameran.
Sex pojkar och två män är bredvid ett stort träd.
En grupp unga män står tillsammans med munnen öppen.
En skallig man med glasögon som bär en grå långärmad tröja och jeans har sin vänstra hand upp mot munnen.
Det finns en man som spelar basket bredvid ett litet barn.
Två barn träffas av en våg i havet
Två leende flickor som håller varandra i handen.
En pojke gör ett trick på sin skateboard i en park.
Grupp av människor som sitter i solstolar på uteplatsen tittar på bergen.
Två äldre kvinnor tar bilder med sin kamera medan en annan äldre kvinna klockor.
Två skidåkare hoppar över en snöhög under starkt solsken.
En kvinna i rosa skjorta rider en häst i en rodeo.
Folk i en parad klädda i mångfärgade kläder och dans.
Tre personer är fåniga i skogen.
Två hockeyspelare slåss med den ena slår den andra i ansiktet.
En kille på en skateboard gör ett stunt i skymningen.
En man i vit skjorta sjunger med ett band.
Snowboardåkaren gör ett trick från sidan av en stor grön byggnad.
Lilla killen i röd snödräkt med hej kattiga vantar
Den här mannen i gul skjorta justerar den blå cykeln för en ung pojke.
En man med lila hatt klättrar på en sten.
En kvinna som försöker sätta på sig ett par strumpbyxor i ett rum utan rum.
En man klättrar upp för en sten.
En person i en blå jacka klättrar upp för en stor sten i en mörk skog.
En pudel som springer längs en strand med en käpp i munnen.
En ung skidåkare får en lektion i snö från en vuxen.
Människor observerar djur i en täckt utställning på zoo.
Människor som går genom en produktionsmarknad med vackra taklampor.
Två män med shorts går upp för trappan.
Två kvinnor med små barn pratar på gatan.
Tre hundar springer mot ett staket i snön.
En man och kvinna och två små barn sitter i golvet med inslagna julklappar.
En vacker vit fågel flyger iväg.
En man i hatt sitter på en soffa med ett spädbarn.
En man med svart hår skär fisk.
En orkester, i formell klänning, med en man som spelar cello i mitten.
En man träffar en volleyboll på stranden.
En liten flicka ler i sin snödräkt medan hon leker i snön.
Två äldre kvinnor som handlar i ett varuhus tittar för närvarande på strumpor.
Den svarta hunden springer genom ett träskigt område med träbitar i munnen.
En man sitter vid en röd byggnad medan han röker.
En kvinna tittar på något som belyses av två glödlampor.
En skara människor som går på gatan med tomten.
Den svarta och bruna hunden jagar något han har sett.
Byggarbetare lägger ut trottoarer för att reparera en väg.
En tjej ska blåsa på en streamer, medan den andra skrattar.
En man som ramlar över i en havsvåg
En basketspelare i svarta hopp, medan en annan i vita försök att blockera.
En liten pojke hoppar upp och ner.
En liten flicka hoppar i balett i klassen som två andra tittar på
Två barn använder beskärningsverktyg på gården.
En svart hund med röd krage springer på snön.
En ensam skateboardåkare som hoppar på en stor skateboardramp.
Ett gäng hundar på en strand.
En man i blått spelar fotboll.
Vissa dansare i kilts tävlar inför en domare i svart.
En kvinna håller ett sovande barn.
En basketspelare har hoppat upp i luften för att skjuta basketbollen.
Den unga kvinnan i blått springer på ett löpband.
En kvinna i topp hatt försöker ta sig in i en maroon bil på natten.
En kvinna applicerar sitt läppstift.
En vit och brun hund, klädd i en bandanna, hoppar genom luften.
Den våta hunden har hämtat den rosa väskan med aqua handtag.
En man som bär en vit tank topp och vit hatt är gravyr nyckelkedjor.
Fem personer sitter på klipporna nära ett träskjul.
Två personer står på en gräsbevuxen bergssluttning framför ett stort träkors.
En svart pudel leker med snön.
En svart pudel springer i snön.
Två gitarrspelare klädda i vitt
En kvinna i baseballhatt och jeans klämmer in en mopp i en gul hink.
En man och kvinnor som äter medan de delar hörlurar.
En grupp elever i uniform lyssnar uppmärksamt på klassens front.
En man står bredvid en BMW.
En liten grupp asiatiska kvinnor samlas under en röd fana.
Två kvinnor på en byggarbetsplats.
En grupp frivilliga hjälper till med att bygga ett hus åt Habitat for Humanity.
Män som jobbar på att bygga ett hus.
En grupp människor som håller i verktyg står framför ett ofullbordat hus.
Fyra arbetare står mellan bjälkarna i ett hus.
Mannen på taket bär solglasögon och arbetar hårt.
En grupp människor utanför med brädor och byggverktyg.
Flera människor bygger en liten byggnad på en fullsatt gård.
Tre tjejer har spikar på ett tak.
Två flickor i en tredje flicka i bymiljö.
Män med kameler samlas på en strand.
Ett blond barn springer nerför sanddynen medan ett annat ser på.
Två hockeyspelare slåss för pucken på hockeymatch.
Tre indiska män sitter tillsammans med korgar med färsk frukt, grönsaker och örter i korgar vid sina fötter.
En man i grön skjorta hoppar i en tvättstuga.
Fyra personer står framför en skåpbil och håller på att bygga.
En man tittar på när en flicka ritar när han äter.
En grupp ungdomar leker med vattenkanoner och står framför en vit lastbil.
En man som knäböjer på ett tak och rör vid en plywoodbit som bär solglasögon.
Man flyger genom luften på skidor över ett berg.
Pojkarna leker med Legos.
En född hund bär lite frukt i munnen medan två andra hundar följer honom.
En skidåkare på ett snöigt skidhopp
En liten flicka sitter på trottoaren och tittar på färgglada barnfärgsböcker.
En mor håller sitt barn på ett tåg.
En man i svart skjorta och tröja tittar ner.
En mountainbikecyklist rider genom en skog.
Någon som cyklar är uppe i luften över en grus- och bergsstig.
Asiatisk kvinna i svarta stövlar och tights med kort klänning lutar igen staket.
En hund är i en del vatten med en trädgren i munnen.
Två afrikaner i röda och blå sjalar poserar för en bild utanför en frisörbutik.
Två barn leker på vägen en snöig dag.
Ett barn sitter på en skidutrustning i snön.
En hund håller en stor käpp i munnen i skogen.
Flickan i skidjackan går nära byggnaderna.
Folk samlas för en bondemarknad dag, handla mat och kläder på en solig dag.
En fågel svävar med vingar breder ut sig.
En pojke står och pekar på en annan pojke som är uppstoppad på golvet.
Två pojkar lade armarna om varandra och poserade.
Två kvinnor är utanför och en kvinna bär ett förkläde som tittar in i en svart maskin.
En kvinna på scenen pekar på en man som håller upp sin hand
En dimsyn av en cykelförare framför en kulle.
En surfare rider många vågor.
En byggnadsarbetare i en orange väst skyfflar stenar medan en annan i en blå väst klockor.
En man med en vit skjorta som håller i ett rack ätbart.
En man med vitt skägg bär ett förkläde och i köket.
Två män spelar i ett band.
En man i vit resaruntskjorta röker bredvid en container.
Dansare poserar framför en flerfärgad, ritad (konst ) bakgrund.
En hund springer längs en strand nära vågorna.
Två små flickor går nerför en stor öken.
En mörkhårig kvinna i svart outfit och svarta höga klackar poserar för en bild med kaktus i bakgrunden.
En liten hund med en boll i munnen som springer genom en kurs.
Två unga pojkar poserar med en person klädd som en Power Ranger.
Folk är på stranden och solar nära klipporna.
Hundarna springer genom vattnet.
En kvinna i roller derby utrustning tittar över rummet.
Mannen är parasailing och gör ett trick.
En grupp människor på skidor med två hundar.
En flicka med blå glasögon och randig baddräkt leker i en simbassäng.
Ett barn som går i snön.
En basebollspelare i blå uniform har precis släppt baseballen på sidlinjen.
Barn som spelar baseball i en allmän park.
Två killar spelar gitarr på scenen med många ljus.
En man tittar upp på en bräda.
Den vita och svarta hunden springer genom ett fält.
Två män i reflekterande kläder som arbetar i en tunnel.
Män som bär ljusgula jackor skjuter gröna bins när andra människor går förbi.
En kvinna som ger en presentation med hjälp av en bildspelsprojektion.
Två män rider en smutscykel och en faller av i en lerpöl.
En säkerhetsvakt står bredvid en ljus orange annons.
En kvinna i en marknadsgester till en hatt, medan ett barn sträcker sig efter hatten.
En tjej i svart och blå våtdräkt surfar.
Den spanske mannen gick mycket snabbt nerför kullen, med sitt barn.
Tre hundar sliter på samma leksak som de står bakom ett hus.
En grupp dansare uppträder under en parad på en stadsgata.
Tre män och två kvinnor som pratar.
Killen låter sin tjej slå honom i ett lokalt cykellopp.
Tre kvinnor står tillsammans och pratar med varandra.
En liten grupp människor chattar på ett torg i staden.
Hunden slickar inuti jordnötssmörburken.
En skateboardare utför ett hopp på en sluttning.
En kvinna som håller ett barn med två barn runt sig
En grupp människor pratar och en annan grupp tittar på fotografier tejpade på väggen.
En svart hund gräver i snön.
En liten flicka med flätor leker med en kamera stativ.
En man är på en skateboard hoppa från en kort avsats på trottoaren.
Två hundar brottas i snön i ett inhägnat område.
Lamm på en gräsbevuxen kulle.
Några kvinnor dansar på en basketmatch på planen.
En man i dagglo gul samlar skräp längs en gata medan andra tittar på.
Person på rullskridskor klädda som clown håller i en skrikande pojke som bär en blå duncehatt och blå trollkarlar cape.
En flicka tittar på ett stativ.
En asiatisk man försöker släcka en löpeld med en liten trähink.
Unga dam målar en annan unga damer ansikte utomhus.
En man fiskar på ett inlopp i havet.
En hund som hoppar för en frisbee i snön.
En kvinna slinker spannmål på marknaden.
Ett litet barn står framför kort vitt bord.
En brun hund i snön har något varmt rosa i munnen.
En man står på en lång plats i en vattenförekomst.
En flintskallig man i en tanktopp som cyklar genom en stad.
En kvinna är utanför en affär och tar en bild och gör ett ansikte.
En person dras av vattenskotrar över det glänsande vattnet.
Två personer och en hund är i snön.
Tre människor, som bär fallskärmar, faller fritt ihop genom himlen.
En brun hund vadar genom vatten och går mot en sten.
En man i svart skjorta tittar på en glaciär.
En man i svart skjorta går på klippor.
En dam sitter på en veranda sving på gården medan en flicka sitter på marken bredvid henne.
En kvinna som bär hjälm rider sin cykel nerför en brant lutning.
En rottweiler bär en mycket lång käpp i munnen genom skogen.
En man sitter i ett gräsbevuxen område och observerar landskapet nedanför.
Ett barn i en Tye-färgad skjorta klättrar på en stenvägg med ett annat barn.
En kvinna håller huvudet mitt i produktionen.
En spansk familj som sitter runt ett bord och njuter av en måltid tillsammans.
Två barn spelar fotboll
En mycket ung leende pojke är i jeans och sneakers står och håller på en bit av gym utrustning utanför.
Tre män sätter saker på sin blå båt.
Den gröna kuperade landsbygden är där folket samlas för att sitta ner.
En äldre man blåser luft i ett föremål.
Den lilla hunden retar den stora hunden på fältet.
En blond man sätter upp ett tält.
Cyklist klädd i svart och vitt med vita solglasögon på poäng på något.
Tjejen i poolen kastar tillbaka håret över huvudet.
En ung kvinna med långt blont hår planterar i en trädgård.
En man i röd skjorta slaktar ett litet djur på en träbräda.
En ung man i baddräkt med vatten som störtar bakom honom.
En brunhårig liten flicka kliar sig i ögat i en barnvagn.
En bred bild av en livlig gata i ett lugn
Ett lyckligt par återvänder från sin shoppingrunda.
Ishockey målvakten är klädd i en röd remsa.
En ung man som stirrar utanför ett restaurangfönster.
En grupp människor som börjar, från startgrinden, på en 5K händelse.
En grupp människor klädde upp sig färgglatt.
En kvinna i grön kostym står framför en topless kvinna med målade bröst.
Folk i en lastbil full av säckar på ett fält fullt av får.
En man hjälper en ung pojke att lära sig att cykla trehjuling.
En snowboardåkare försöker hoppa på en pysselåkare.
En kvinna i svart jacka och en man i vit skjorta passerar varandra på trottoaren.
En hockey målvakt hukar på isen.
En pojke med blå skjorta går nerför en rutschkana.
En kvinna som vandrar i snön med hjälp av skidstavar.
Killen i den vita uniformen har en basketboll i handen.
En basketspelare dribblar bollen under en match.
En person som gör ett cykelhopp, en skyline i bakgrunden.
Två män pratar medan en till tittar på.
Damen håller sin pensel bredvid konstnärens staffli.
En kvinna med vit skjorta går på trottoaren med en stor sopare.
Två män hoppar upp för bollen nära bågen i en basketmatch.
En kvinna i röd rock är på skidåkningen.
En kvinna i svart hatt pratar med en kvinna i blå klänning.
En kvinna i blå skjorta och halmhatt målar utomhus.
Folk går nerför gatan och förbi en öppen buss.
Grupp av män och kvinnor som väntar på en buss.
Flera män klädda i bakoveraller sjunger och spelar instrument.
En hockeyspelare ser kraftigt nedåt.
En person rider en skateboard i luften ovanför en ramp.
Tre män med gula arbetsvästar står bland en grupp människor.
En kvinna i röd jacka och en annan person får ut sina snowboards på en snöfylld parkeringsplats.
Kvinnan svepte en flagga runt sin kropp och brände rökelse.
Ett par går nerför en livlig stadsgata när de passerar en fågelshow.
En kvinna och två manliga musiker med musikutrustning.
En man på maskinen pratar med en kille klädd i en galen utstyrsel.
En kvinna som håller i en klädkorg framför en byggnad med en lägenhet att hyra.
Pojken i blått har bollen, och pojken i vitt är luftburen.
En man glider en skateboard nerför en trappa ramp.
Två äldre kvinnor sitter på en träbänk utomhus.
Två hundar jagar ett klippt gräsfält.
En person cyklar på en stig bredvid skogen.
En mor och hennes tre barn går på en gata.
Tre honor och en hane går vid kanten av en väg.
Den bruna och svarta hunden springer över gräset.
Två barn står i gräset och sprejas av en slang.
En rödklädd man spelar gitarr på gräset.
En grupp barn som bär blå och gula uniformer sätter ihop händerna.
En dirt bike rider är i luften drar av ett trick.
Två asiatiska flickor klädda i svart poserar för en bild framför torra träd.
En ung vuxen dansar på sin hand.
En snowboardåkare med grön jacka hoppar över en låg grind.
Ungdomar övar på att gå på den höga tråden.
Pojke med blå huva hoppar över ett trappräcke.
Två asiatiska flickor sitter på ett blomsterfält.
En skateboardåkare är i luften efter att ha åkt upp för en cementramp.
En skidåkare som slingrar sig nerför en bergsstig.
Två unga flickor rider beige camels som en annan dam bär en handväska klockor.
Två honor rider kameler baklänges.
En man i orange är böjd över att svetsa något på marken.
Två personer i skyddande redskapssvetsning.
En grupp pojkar leker på en strand.
Ett gathörn med parkerade bilar - vita, röda och tillbaka.
En man med glasögon stirrar på kameran.
En flicka hukar sig på en skateboard bredvid en färgglad vägg.
En välbalanserad hane står på ena foten nära ett rent havsstrandsområde.
Två unga flickor pratar med en man i en skåpbil.
Pojkarna spelar fotboll på deras kvartersgata.
En liten asiatisk flicka äter snacks medan hon ler mjukt.
En liten grupp människor som observerar vildmarken under dagtid.
Tre personer på gör högriskjobb.
Många människor är utspridda längs en strand eller lagun roar sig.
Två unga älskare som håller på att gå skilda vägar.
En grupp människor sitter under ett plåttak.
Vänner som skrattar åt något de just har bevittnat.
Många människor går i staden nära höga byggnader.
En man Rollerblades på en skridskobana.
En grupp afrikanska kvinnor och barn som bär färggranna kläder.
En grupp barn som sitter mot en stor röd container.
En kvinna som fotograferar ett föremål på en säng.
En pojke på en svart surfbräda rider vågen på magen.
En klättrare med gul ryggsäck går längs åsen på en snöig bergssluttning.
Två män spelar gitarr tillsammans
En person på en snowboard hoppar över en klippa i snön.
En afrikansk kvinna står med sina två barn under ett stenblock.
En man och ett barn pratar en promenad genom en park.
En man ger en låda till en annan man i en grupp.
En grupp män väntar i kön för att få mat vid ett fönster.
En vandrare går uppför berget på en snötäckt väg.
En ung pojke hoppar upp i luften med hjälp av en studsmatta.
En flicka och en kvinna rider en kamel.
En cowgirl lassoar en ung vit kalv från baksidan av sin bruna häst.
Två blonda kvinnliga brottare i ringen.
Kvinnan i den röda jackan tittar på barnet i en grön jacka.
En man och en kvinna visar sina tatuerade hjärtan på sina handleder
Två personer står på tre hästar som en del av en parad.
Vissa människor väntar på att korsa en livlig gata i Portland Oregon.
Indiska studenter arbetar och diskuterar i ett klassrum.
Ett barn håller tre fåglar i sina händer.
Skidåkare hoppar högt framför träd i snöigt vinterlandskap.
En gul motorcykel kör nerför vägen.
En person observerar bilder som är i ramar på en vägg.
En man på en motorcykel kastar en wheelie i smutsen.
Afrikanska barn i en brunn med en hämta vatten genom att dra upp en hink.
En brun och vit hund bar tänderna i snön.
En afrikansk familj samlades utanför och förberedde något i en gryta över en eldsvåda.
En grupp människor springer nerför en gata.
En restaurangs bås är ljust upplysta och omgivna av speglar.
En skidåkare som bär blå snöbyxa flyger genom luften nära ett hopp.
En speciell dagtavla på en restaurang.
Två hockeylag tävlar.
Många människor går längs en stig bredvid en lång byggnad och träd.
En vit hund med svart krage springer i snön.
En man raderar en liten dunge lastad med gröna växter på en flod.
Några kvinnor och barn är på trottoaren.
En kvinna pratar med en man som håller i ett glas öl.
En ensam skidåkare som åker genom snön.
En tonårspojke rider på en skateboard utanför en tegelbyggnad.
En stuntcyklist hoppar upp i luften bredvid den nedgående solen.
En man på en cykel i luften
En vit hund har fångat en pinne på stranden vid havet.
Tre män och en liten pojke jobbar på ett grönt modelltåg utanför.
En kvinna i svart konverserande går längs trottoaren en kall dag.
En asiatisk flicka står i folkmassan och bär rött läppstift.
Ensamhetsbåten flyter på sjön.
Två hundar är på en stig i skogen medan två människor tittar på dem bakifrån.
Barn spelar monopol tillsammans.
Tre kvinnor i amerikansk kolonialstil sitter tillsammans och syr.
En ung asiatisk flicka står mellan två trädstammar.
Tre ryttare bär svarta tröjor hoppar sina BMX cyklar i luften.
En konstnär som skulpterar sin staty.
En gammal kvinna har påsar på en livlig gata.
En hund som leker boll i sanden.
En man i ränder och en i läder poserar för kameran i en stad.
Två gamla män i vinterrock går genom skogen.
En man på en buss som tittar framåt.
Två personer går förbi ett gammalt hus.
En snowboardåkare gör ett stort hopp och är i luften.
En mur med skrifter från arga demonstranter i en stor stad.
Det finns 5 bruna hundar på koppel med sina ägare i närheten.
Tre vita hundar är nära en svart lama.
En man i smoking spelar ett mässingsinstrument i ackompanjemang med en kvinnlig pianospelare.
En blond tjej läser pojkscouthandboken.
En stor brun och vit hund hoppar genom håret.
En parad av inbördeskrigssoldater som spelar flöjter och trummor.
En grupp killar som spelar basket i en park.
Två kvinnor böjer sig över för att röra vid en liten känguru.
En kvinna ligger i en säng med blommor på filten.
En glad man slår läger ute i snön med rosa flamingos.
En man med solglasögon sitter på ett däck.
En grupp hundar leker tillsammans i snö.
En grupp människor står framför en försäljares monter.
En grupp män hejar med styrofaamkoppar.
En orientalisk kvinna tittar på en liten uppvisning av kosmetika på ett bord.
En ung flicka har en grön plastlapp, tjejen i lila är i köket bakom henne.
En man med glasögon och skjorta som säger "fick stenar?" vänder en pannkaka ur en stekpanna.
En grupp människor som tittar på en snowboardåkare utför ett trick.
Personen i den svarta skjortan utförde ett stunt på gatan medan publiken tittade.
En fallskärmsåkare lyfter från marken.
En grupp människor står framför vissa butiker.
Två killar är i ett gym, den ena tittar på den andra träffade en tung väska.
En man och en ung pojke sitter på ett steg och äter apelsiner.
Tre dansare med röda stygn uppträder på en mörk scen.
En grupp människor tittar på färsk sallad på den lokala gatumarknaden.
Flera personer står utanför och sjunger i blå och gröna kläder.
Unge pojke i vit baddräkt hoppar upp i poolen.
Den unga dansaren marscherar i paraden.
En pojke på en skateboard som glider på en räls.
Två BMX-cyklister på en lerig kurs.
En man i rött och svart slår en fotboll med huvudet.
En stor fågel flaxar sina vingar över vattnet.
En hund springer över snön med en stor käpp i munnen.
Baseball spelare bär guld hjälm med blå jersey och grå byxor.
En utfältare som är på väg att fånga en flugboll.
Två baseballspelare byter handslag.
En vit och brun hund springer uppför en gräsbevuxen kulle.
En kvinna köper en stor mängd kattskräp från en Walmartbutik.
En man i jeans och en grön skjorta jobbar på en hockeyrink.
Ett litet barn skriker med människor omkring sig.
En cykelförare tar ett djärvt hopp när hans vänner tittar på.
En brun hund springer på brunt gräs.
En basebollspelare i en blå uniform slår en löpare till basen.
En baseballspelare springer till basen.
En man kastar en boll över fältet.
Mannen i den röda skjortan bär en svart väska genom stadens gator.
En äldre asiatisk man bär en svart och grön jacka och en New York-hatt med cykeluthyrningsskylt.
Två kvinnor i svart tränar kasta gevär i luften.
En svart hund hoppar ner i vattnet och fångar en käpp i munnen.
En gammal asiatisk man i röd mössa och blå jacka ler.
En skara ungdomar dansar i mörkret.
Ett skolband går i en parad.
Den här stora svarta och vita hunden springer på sanden.
En tjurryttare har precis flugit från en häst.
Utsikt över en fotbollsboll sparkas in i ett målnät
Två små flickor sitter på en lejonstaty.
Två pojkar paddlar över vattnet med fiskenät, den ena bär en långärmad gul skjorta och den andra bär en påse hoodie.
En man åker nedförsbacke på ett berg.
En kvinna med mörkt lockigt hår och en mörk klänning sjunger och håller i en gitarr.
En underbar dam som spelar musik.
En kvinna med svart hår med lila ränder i det tar ett bett medan hennes följeslagare i en röd skjorta ser på.
En brun hund som springer genom det smutsiga leriga gräset
En man som bär en sportuniform går nerför fältet när en annan följer efter.
En medelålders man som vilar efter trapetsen på cirkusen.
En kvinna i svart skjorta stoppar en sked i munnen.
En liten flicka som rider på en leksakshäst under julen.
Två kvinnor som bär vita badrockar slappnar av på en soffa med fötterna uppsparkade på ett soffbord.
Folk som dansar framför instruktören
Två kvinnor i baddräkt leker på stranden.
Två kvinnor sitter på en skidlift, med berg i bakgrunden.
En ung pojke klänger sig fast vid benet på marmorstatyn av en barbröstad kvinna.
En asiatisk kvinna i svart bikini tittar på en mobiltelefon nära poolen.
En svart och brun hund brottas, och en liten hund klockor.
En blond kvinna gissar på en brunhårig man på kinden.
En orkester som övar och spelar musik i en sal utan publik.
En man som står i en vit skjorta leder en liten grupp violinspelare.
Någon går genom snön med snötäckta berg bakom sig.
Människor med utrustning klättrar upp för ett snöigt berg
En pojke med mörk och en kvinna i brun skjorta leker med en lila uppstoppad leksak.
En liten flicka som klättrar på en repapparat.
Två män går längs en livlig stadsgata med ord tryckta på trottoaren.
En man i en mörkfärgad tröja och står bakom en stol.
En grupp människor står ljud utomhus, en bär rosa byxor och en blå topp.
En Notre Dame baseballspelare som sköter baserna.
Två killar är på ett baseballfält och en är på väg att träffa basen.a grupp
En grupp människor som sitter på avstånd.
Med höga glittrande vita kronor poserar en man och en kvinna tillsammans med palmstress och glittrande röda och vita stjärnor i bakgrunden.
En man står på en häst framför en publik.
En person som bär klänning går längs vattnet i leran.
En arbetare reparerar tegel på en skorsten.
Skateboarder på en ramp som syns genom ett kedjelänkstaket.
Person som sitter vid ett skrivbord i ett bibliotek.
En baseballspelare försöker glida in i tredje basen medan en annan spelare blockerar honom, när en umpire närmar sig.
En baseballspelare i vitt svänger på bollen.
En kanna gör sig redo att kasta en boll under en basebollmatch.
En av spelarna spelar för det irländska laget.
Att försöka hålla fast är lika mycket en bra idé som en dålig!
Mannen fyller sin bil med bensin.
En man använder en patron rakhyvel för att raka kinden.
Fem gamla män som spelar pool
Två kvinnor går framför en buss för att korsa vägen.
En röd bogserbåt ska docka i en hamn.
En hund hoppar i luften parallellt med en tennisboll.
Två barn kör över en sanddyn.
En kvinna hoppar på toppen av en sandkulle.
Tjejer deltar i en basketmatch framför en publik.
Arbetare skapar ett föremål av metall och trä.
Tjej i rutig skjorta som rider enhjuling.
Tre män går i rad, den ena bakom den andra, på en gata framför en affär som heter "The Odeon".
En grupp vänner glider nerför en sandig kulle.
En längdskidare grimaserar när han klättrar en liten lutning.
En man i hatt som sover i en stor brun stol.
En liten flicka i klargrön går på trottoaren medan hon bär en väska eller låda.
Två män väntar på att bli intervjuade, medan en annan kollar mikrofonerna.
En kvinna scoopar glass medan en man sitter vid bordet bredvid henne.
En kvinna med långt brunt hår sitter ensam i en bar.
En liten blond flicka i grön parka och röda regnstövlar placerar en fot vid kanten av en liten sjö, med vintriga träd och en ockuperad utombordare motorbåt i bakgrunden.
Två skäggiga män och en kvinna.
En folkmassa full av människor håller flaggor och skyltar.
Fyra barn klättrar uppför en snöig kulle, en kämpar.
Två män i en gränd, en med händerna i fickorna och tittar åt ett håll bakom honom.
Tolv personer är redo att lyfta i en varmluftsballong.
En man sitter på en bänk nära stranden och knyter sin sko.
En man spelar gitarr på trottoaren.
Två män Nordic ski racing medan andra tittar bakifrån.
En grupp på tjugo män sitter runt ett bord.
En person åker skridskor längs insidan av ett långt rör.
En surfare rider på en våg.
En man cyklar genom ett skogsområde på morgonen.
Folk på trottoaren, medan en person på gatan håller en yxa.
En pojke är luftburen på en cykel ovanför en stadspromenad nära en ledstång.
Muzzled greyhounds tävlar längs en hundbana.
En man med långa ärmar skjuter på natten.
En rödhårig kvinna med folk i bakgrunden.
Tre hundar ligger i snön framför ett stängsel.
En person som sitter på en hiss över vatten med en annan person lämnar en väska till dem.
Pojken sitter på en soffa och stirrar med en hammare i händerna.
Snowboardåkare gör tricks på berget.
En person på en motorcykel som gör en wheelie från en sten.
Flickan i den gula klänningen ser så söt ut.
En pojke och hans hund står på en studsmatta och njuter av varandras sällskap.
En ung kvinna som tvättar sin bil.
En man håller och tittar på en produkt i en livsmedelsbutik.
En fågel, vingar över vattnet.
En liten flicka i gul klänning sitter på de vita klipporna.
Ett barn gör sig redo att glida ner för rutschkanan.
En kvinna i en affär håller ett föremål i sin vänstra hand medan hon tittar bort från kameran.
En person hoppar en cykel från en ramp i en karg skog.
Två unga kvinnor ska korsa gatan när en gul skolbuss passerar.
En äldre kvinna bär en rosa randig skjorta.
Man sitter i en svart stol och röker på en restaurang.
Folk slappnar av i gräset på natten under en karneval.
En kvinna i svart och orange jacka kastar en pinne för en brun och svart hund att hämta.
En stor grå och vit vattenfågel.
Två hundar leker med varandra på gräset.
Folk rider på stranden.
Folk i orange rock ställer sig bakom en man som bär solglasögon.
En manlig skateboardåkare drar nytta av halvröret.
Den grå och vita hunden springer genom snön.
En grupp tjejer äter ute på däck.
En grupp vänner leker i en sjö.
Surfaren passerar en annan surfare medan han paddlar in i surfingen.
En kvinna på sin laptop ler mot en person i en blå skjorta bredvid henne.
En kvinna i laxfärgad skjorta talar och ger gester till en man i grön skjorta.
En man parkerar sin cykel utanför en byggnad bredvid en staty av en mans huvud.
En kvinna i brun skjorta som pratar på en rosa mobil.
En person i en regnrock står i en båt som går över vattnet.
Skidåkare i rött hoppande högt i luften över snön.
Liten brun hund sticker huvudet i en coloful väska fylld med tyg.
En flicka glider in i basen under en softball spel.
En person städar upp en röra framför en scen.
En grupp människor är i vattnet.
Fem män som bär smoking hoppar upp i luften framför en liten flod
Mannen och hans två barn är på väg att gå förbi en person.
Två hundar skäller i ett kök medan en person sitter vid ett bord.
Den här personen fallskärmshoppar med skidor upp på en snöig kulle.
Två män och två kvinnor i jackor går nerför en stor stad gata.
Två kvinnor pratar med varandra utanför.
En man är i luften upp och ner i snön.
En man tittar på konstverk.
En hund är på toppen av en blå bild och en liten pojke är bakom honom.
En softball spelare försöker desperat att nå sin bas medan motståndaren taggar ut henne.
Två kvinnor med långt hår och storbonade fysiker poserar för en kamera framför träd.
Ett par män som sitter utanför en bar
En person i en rutig skjorta tar en bild av en vit vespapåse på något gräs.
Ett litet barn leker på en strand bredvid en tom stol.
Folk står i en byggnad som är under uppbyggnad nära 3rd St.
En pojke och hans husdjur padda bara umgås.
En man som bär en ha tar sin häst ut på en promenad.
Folk äter ute på ett väldigt långt bord.
En man i blå overall hänger från en metallstolpe med en sele.
En liten grupp människor tittar på en konstnärlig vattenfontän.
En person som sitter i en grön stol utanför en byggnad omgiven av skräp.
En vit man med blont hår dricker öl.
Ett lag fotbollspelare lyfter en lagkamrat så att han kan nå bollen.
Mannen med spetsigt hår sitter vid en färgglad affisch.
En gammal man håller i kopplet på en vit mula som drar en röd kärra.
En snowboardåkare tar sin bräda när han är i luften.
En pojke står på en snöig kulle och tittar på en solnedgång eller soluppgång.
En liten hund jagar en vit boll på gräset
En person som bär kinesisk hatt, trädgårdsskötsel, medan en grupp människor som står i motsatt riktning står bakom honom.
Skateboardåkaren vänder sig om och håller sig på marken.
En man i röd tröja håller ett barn ovanpå axlarna.
En blondhårig liten pojke som klipper sig.
Ett barn med cowboyhatt sitter med gitarr i knät.
En liten babyklänning i gula leenden.
Flickan pekar på en gejser
Två hundar springer över skogen.
En person med livliga kläder som dansar på lite betong.
En snowboardåkare hoppar över en tunna.
En man klädd i vitt med en vit mask i ansiktet som låtsas vara en staty på en plaza.
En man i krageskjorta håller en babyhand.
En man och hans barn tar en bild med kuddar över huvudet.
En blöt hund stänker genom vattnet.
En man som hoppar med en skateboard under en bro.
Folk går framför Outdoor World-butiken.
Kvinnan i blått verkar blåsa glas medan ett barn tittar på.
Pojken i flerfärgad randig skjorta tittar på den röda lådan.
En ung man som bär kostym, slips och solglasögon går nerför en trottoar och håller upp ett papper i läsningsstil.
Den stora bruna hunden satt på sängen överväldigad av omslagspapper.
En man använder en maskin på marken framför en sten påfågel.
Hunden simmar och plaskar genom vattnet.
En liten pojke tittar på en liten flicka i vitt cykla med träd.
En hund slickar näsan.
En svart och brun hund som leker med en pinne
En man i jeans som håller en cykelram med en annan man i bakgrunden.
Man med orange duffel väska och flicka i grissvans knuffar en laddad vagn ner för en trottoar.
En hund hoppar över en bar med en boll i munnen.
En kran, vingarna över havet.
Hunden vilar efter en omgång hämtning.
Ett leende litet barn sitter i ett badkar med sitt våta hår draget i en lång, våt spik som kommer från toppen av hennes huvud.
En skidåkare som gör ett trick på stången medan han fotograferas av en annan man
Två bruna hundar slåss lekfullt i snön.
Två kvinnor hjälper en brud med sin bröllopsklänning.
Ett par barn som är utanför, försöker på inbördeskrig era kläder.
En man åker snowboard nerför en snöig kulle.
En man sitter på en cykel mitt i skogen.
En man cyklar på en kulle.
Hane med vit skjorta och brun jacka som sitter bredvid en hög bönor.
En muslimsk man som bär solglasögon lagar mat.
En snowboardåkare som bär en röd jacka går nerför ett berg.
En flicka lockar i en tävling.
Tre tonårspojkar i t-shirts går nerför gatan.
En man som städar vid fönsterglaset
En ung man lyfter en stor skivstång i ett gym.
Två män jobbar på en bogserbåt.
En kvinnlig sångare klädd i en solbränd klänning drar en mikrofon mot henne när tre musiker som spelar stränginstrument ger musiken.
Det är en person som spelar gitarr.
En mamma som håller sitt barn i knät.
En kvinna i en vit outfut spelar tennis.
I ett tomt fitnesscenter hukar sig en kvinna och förbereder sig för att lyfta en lång vikt.
Många bestämmer sig för att det är dags att äta.
Två kvinnor i svart har blod på ansikte och knä.
En brun hund springer längs gräset.
Två unga asiater, en flicka och en pojke, klädda i kostym, sitter vid ett bord och tycks studera.
En bild på Jim som bär glasögon i en labbrock.
Två män skiner sina kunders skor utanför.
Två lag tävlar i en fotbollsmatch.
Fiskare vid sandstranden sida vid sida kastar nätet till havet.
Den här mannen är på en restaurang som har spelautomater.
En man i vitt och grönt spelar fotboll på ett plan.
Två flickor i blå uniformer en tjej i vitt spelar fotboll.
Två figurer står i en snöig miljö klädd i vita och varma rosa kläder, stirrar mot ett berg.
Folk tittar på flygplan i en stor händelse.
En orientalisk kvinna som bär svart tunika, leggings och stövlar står utanför en produktaffär.
En cyklist flyger genom luften nära sanddyner.
Ett par tittar i vördnad på en utställning på en karneval
En hund fångar en leksak i snön.
En liten flicka drar på en filt medan en liten pojke ligger ovanpå den.
Två flickor som spelar i en park.
Tre unga studenter sitter vid bord i biblioteket och arbetar med läxor.
En ung pojke hoppar från en klippa i skogen
Den svarta och vita hunden hoppar vid en stock nära en bäck.
Man och kvinna på natten dansar med snurrande facklor i händerna.
En man i glasögon sitter bakom ett bord fyllt med militära minnesmärken.
Brun och vit hund som rullar runt på gräset.
En kvinna i brun väst går på snön med ett djur.
Det finns en hund som springer längs stranden.
En man i solglasögon, en röd randig tröja och en skinnjacka ler och pekar finger.
Två män jobbar på Apple laptops.
Blöt brun hund, hoppar upp ur vattnet.
En uniformerad man tittar på tåghastigheten.
Två arbetare med gula hattar och blå arbetskläder städar en parkeringsplats.
En man i mörka kläder lutar sig mot en byggnadsingång med upphöjda armar.
En pojke på en skateboard som maler ner en ledstång.
En basketspelare kör till korgen.
En manlig basketspelare håller fast vid kanten av ett basketmål.
Två lag som spelar rugby i marken.
En fotbollsspelare i rött blir träffad av en spelare i vitt.
Två kvinnliga fotbollsspelare tävlar i ett spel.
Mannen till vänster tittar på kvinnan och mannen.
Tre små barn som rider på en åsna dragen vagn.
En man som bär svart skjorta och glasögon höjer händerna medan han sitter vid ett pokerbord.
Två basketspelare på motsatta lag längtar efter bollen.
En basketbollspelare kommer ner efter att ha doppat bollen.
Många människor bevittnar en fotbollsspelare fånga bollen
En fotbollsspelare i en grön och guld uniform vaggar bollen när han hoppar över en motsatt spelare.
Unga kvinnor spelar ett intensivt spel av lacrosse.
En lacrossespelare firar med en lagkamrat.
Ett litet barn svänger tillbaka mycket högt.
Folk i en skola cafeteria med en pojke i förgrunden bär gula och bruna ränder
Två unga kvinnor poserar och håller varandra i närbild.
En brun och vit hund på studsmatta med skog i bakgrunden.
En man med svart hatt står och skuggar ögonen.
En person som bär grå jacka och solglasögon poserar för kameran.
Två kvinnor med barnvagn i en tjusig restaurang.
En kampsportskonstnär får ett slag mot sin motståndares lår medan en domare kastar upp handen.
En man i en tröja spelar dart.
En grupp säckpipare går nerför en gata i en parad.
Person med skidor och hund står i snön.
En man på en gul surfbräda rider en lätt våg.
Två personer som jobbar på en stege för att få något från ett träd.
En pojke på en skateboard rider på en stenvägg
En cyklist rider på ramper.
En kvinna i mörk skjorta och glasögon tittar på en digitalkamera.
Två män som är i en match med varandra.
Två killar, båda bär vita kostymer en med svart bälte den andra med svart och rött bälte, de har en match.
Mannen i gul kajak paddlar genom forsarna.
En hund som leker i snön med en vit boll.
En kvinna i rosa skjorta tittar på vattnet.
Dansaren får sin sista makeup innan hon går ut på scenen.
Äldre man i rullstol tigger om allmosor
En person springer vid vattenbrynet vid havet.
En man uppträder på stranden.
En grupp vänner spelar instrument mitt i skogen.
En man sover på en bänk utanför.
Folk på gatan kantade med höga solbrända byggnader.
En vuxen ler med ett barn på en gunga.
En svart hund slåss med en brun hund i snön.
En man som bär en fluga och glasögon poserar för ett foto.
Två unga män står med en skylt mot en vägg.
En person som klär sig i svart sitter på en bro.
Två kvinnor med armarna om varandra ler in i kameran.
En man som håller i en drink poserar med en kvinna.
En man kastar en liten vit boll mot några röda koppar.
En man och en kvinna är avslappnade på soffan.
En asiatisk pojke och flicka som går bland en folkmassa med träd över sin stig.
Man spelar en brun och vit elgitarr.
En tennisspelare som gör sig redo att backhand bollen i en tennismatch.
En svart hund hoppar nerför en snöig kulle.
En grupp människor med handskar på arbete på stora färgglada rutor.
En familj som sitter framför ett gräddhus på trappan.
Fem unga män uppträder bredvid ett fönster.
Fem personer är ute i ett parkliknande område och en av dem sträcker sig efter en handsving.
En ensam demonstranter i en svart jacka på trottoaren.
Folk sitter på stolar med utsikt över en brant stenig lutning.
En person hoppar över ett hus på skidor.
Detta är en liten stämpel med blå himmel och vita linjer med gröna buskar.
En brun hund som gräver ett hål framför en växt
En liten pojke på en grön släde på natten.
En stor brun hund skakar av sig i vattnet.
En våt hund kommer fram ur djupt vatten.
En grupp unga pojkar i blå baddräkter försöker hoppa in i en pool till sina simlärare.
En paraskier landar på ett berg.
En kvinna sorterar saker på en ljusblå duk.
En ung man som rullar upp ärmarna på tröjan.
En man använder en lövblåsare för att få löv från trottoaren
En kvinna med en röd baskettröja håller en basketboll och tittar upp.
Två kvinnor sitter vid skrivbord i ett stort rum med vita väggar.
En pojke som håller en läskburk i ett vattenfall
En surfare rider en våg i en stor vattenförekomst.
En ensam man går på en kyrkogård.
En vit hund i en flod jagar en anka
En hund med orange jacka ligger i snön
En grupp asiatiska flickor klädda i rosa och lila poserar i en rak linje
En person i skyddsutrustning som kör en smutscykel.
En man på en släde dras genom snön av sina hundar.
Rödhårig flicka på bakgården som sitter på en såg.
En grupp människor sitter utanför en restaurang i en skidstuga.
Tre män med gröna t-shirts gör en gatuföreställning.
En stor grå fågel med gula ben flyger nära vattnet.
En tjej i rosa leende för kameran.
En flicka i rosa strumpor som hoppar med händerna i luften.
En kvinna håller en kokosnöt framför en intresserad hund.
En ung pojke i randig tröja och jeans som springer i gräset.
En man sitter på en bänk med några väskor.
Under en ishockeymatch försöker en man göra ett mål.
Tjejer i kostymer står och ler.
Två hundar springer genom smuts och ogräs.
En hund går genom snön.
En svart och vit hund springer över ett snötäckt fält.
En hund hoppar genom vatten.
Två unga kvinnor som pratar vid ett bord på ett café.
Ett par kysser varandra på en bro.
En kille som åker snowboard på en sluttning.
Ett litet barn som jagar en pidgin.
En svart och en brun hund går genom skogen.
Två kvinnor sitter vid ett bord med tomma glasögon framför sig.
En hund med en käpp i munnen springer i en skog.
En danstrupp av afroamerikanska ungdomar som gör ett koreograferat drag.
En rad fåglar sitter framför ett grått moln.
Någon tittar på den vackra utsikten över staden.
En man i mitten av avdelningen för kvinnors livsstilstidningar läser en tidning som förklarar "Jag är gravid!"
En svart limousin står parkerad bredvid en trång trappa.
En dam som bär en slaktares förkläde sjunger på en scen medan hennes band spelar bakom henne
En barfota kille i orange skjorta och svarta byxor som hoppar på en studsmatta i en bur.
Ett gäng hundar tävlar i en tävling.
En karneval mitt på natten.
En man i grön skjorta ligger på gräset med en bandanna över ögonen, bredvid en svart fågel.
En kille kör en trehjulig motorcykel.
Ett barn uppträder med en leksak medan på scenen med en färgglad ballong bakgrund.
En grupp människor som går tvärs över en gata
En grupp barn pratar med en tjänsteman.
En man med en röd spansk skjorta och en kvinna med lila ränder i håret.
En cyklist går nerför en grusväg i skogen.
En hund hoppar ur en bäck.
Flera barn i kläder är i ett mörkt rum, och två av dem håller i rep i luften.
En flicka med lila skjorta och solbrända shorts är poserad i ett dansdrag.
En vit hund försöker fånga en tennisboll högt i luften.
En leende man med hörlurar och grå mustasch
En liten blond flicka är insvept i en Care Bears filt med julpapper bakom sig.
En pelikandykning mot vattnet med fötterna ut.
En tonårspojke gör tricks på sin skateboard i ett område med mycket graffiti.
En man som paddlar forsar.
En asiatisk kvinnlig tennisspelare förbereder sig för återkomst av volley på en hälsning och lila court.
En man i flera färger som rider på en surfbräda på en våg.
Ett barn sitter på en trottoarkant med inline skridskor och skyddsutrustning.
Människorna i den röda parasailen glider över vattnet.
En man rider på en bräda i havet och dras uppifrån.
En flicka som utför en rytmisk gymnastik rutin.
Tunnelbanearbetare använder stegar för att kolla in ett möjligt problem som en röd tunnelbanebil flyger förbi.
Fiskare bär poncho och hatt sitter vid kanten av vattnet.
En hund står upp mot armbågarna i snö.
Tre personer står på en stig genom skogen.
En snowboardåkare vänder upp och ner med en snötäckt backe i bakgrunden.
Två kvinnliga gymnast jobbar upp innan deras tur är uppe.
En pojke läser en serietidning framför en röd stol och en grill.
Smutscyklist gör sig redo att börja nedför sluttningen.
Killar som bär gult, rött och blått springer i gräset.
En man i brun väst och glasögon leker med en brun hund.
En flicka i klänning går medan en familj står i bakgrunden.
En ung pojke som försöker spela hacky säck.
Två flickor hoppar högt framför tallarna.
Gamle man som lär lille unge att köra.
En ung kvinna i en svart tank-top tittar och flyr från något bakom henne.
Ett litet barn som sitter i en enda röra av färg.
Två hundar leker och rullar runt med varandra i gräset.
En man som rider en tjur på en rodeo.
Barnen leker i sanden omgiven av en sandstruktur med en hel del fönster som öppningar.
En kvinna på en cykel stannar för att prata med en gentleman som sitter på en stol på trottoaren.
En hund springer med en annan hund i bakgrunden och håller en boll i munnen.
En parad av säckpipare går genom en stad gata.
En ridhäst är på en häst som hoppar över ett plan som ligger på marken.
En man visar upp sitt exibit för många människor.
Den här mannen, som bär ett blått pannband och vit skjorta, spelar tennis.
Två män i solglasögon sitter vid ett bord och dricker öl.
En hund springer i snön och bär på en röd frisbee.
Flera musiker spelar vid en formell social sammankomst tillsammans med två dansare som uppträder.
En man och pojke letar efter något på marken.
Barn och vuxna i ljusa kläder dansar.
En ung dalmatier bär hatt bredvid ett träd.
En dam i en rutig klänning smeker sin vita hunds ansikte.
En pojke jobbar på ett projekt i butiksklassen.
Mannen med blå jeansshorts grillar.
En lacrosse spelare tittar på ett objekt i himlen som inte är bollen.
En grupp unga pojkar leker lacrosse utanför.
En kvinna och en ung flicka sitter ner och ler.
En vuxen man bär en outfit gjord av en Spider-Man sängöverkast.
En tjej i huvtröja tar en tupplur med sin svarta hund.
Skateboarder i grön skjorta gör tricks i luften.
Tre barn i en by står under en markis
En man med en blå väska lämnar en stadsbuss.
Fyra personer, två i gröna uniformer och två i röda uniformer, spelar ett spel av lacrosse.
En man i blå skjorta snurrar en lerskål.
En man i en ljusblå skjorta med en gul och svart halsduk gör en lerplatta.
En man i en röd tröja skjuter upp ett jättelikt träd i en snöig skog.
En ung man i svart och vit randig skjorta vilar på gräset medan trafiken passerar i närheten på vägen.
Två honor med glasögon som går i street arm i arm.
Två små barn står bredvid en fönstervisning.
En massa människor tittar på ett barn i badkaret.
En man sitter på en bänk framför en övergiven byggnad.
En brud som har en fotografering utomhus runt massor av människor.
Golfare i en vit mössa sätta i ett hål medan omgiven av åskådare och andra golfare.
En svart hund som springer i gräs.
En gul hund springer på ett fält nära ett berg.
En mörkbrun hund som står på byggutrustning.
En tennisspelare gör sig redo att lämna tillbaka bollen.
Tennisspelare gör sig redo att spela tennis.
En man med vit hatt svänger armen tillbaka för att kasta.
En man svingar sin klubb i en golfmatch.
En man i en röd kajak trampar genom en våg
Man föreläser för intresserade människor framför en nyckelstaty.
Två män och en kvinna som skjuter på en bar.
Ett par som bor tillsammans med sina barn och blir döpta av en präst.
En man i hatt och jacka står på trottoaren med en hög med skräp framför sig.
Män sitter utomhus under ett träd i full blom.
Folk i köket på en fest med mat och dryck.
Två små flickor som spelar i en flerfärgad bollpenna.
En tonåring i randiga shorts hoppar upp i luften på stranden.
Kayak rider höjer armarna när han är stänkt med vatten.
En svart man applåderar en löpare i röd tröja och nummer 281.
En stor grupp människor tittar på en person som klättrar på en stolpe.
En man i blå skjorta lyfter upp sin tennisracket och ler.
En tonårspojke som gör ett cykeltrick på en cykelramp
Pojken står på lekplatsutrustningen i den blå triangeln.
En man som kysser en pojke i en skåpbil.
Ett barn visar två leksaker medan det sitter i en VW-buss.
Två blå uppblåsbara flottar är inblandade i en kollision på vitt vatten.
En ljusbrun hund hoppar över ett hinder inomhus.
En individ åker skidor nerför en bergssluttning.
En bäver på stranden av en bäck.
Serena Williams slår en boll i en orange utstyrsel
Två löpare som bär tävlingslappar klättrar över ett träd som ligger tvärs över stigen.
En kille och en tjej som leker med varandra när de sitter på stolar.
Man i brunt och rött rutig knapp upp skjorta och blå jeans gör en manlig och kvinnlig skratt.
Ett barn som springer genom ett fält av gula blommor.
Vissa människor står i ett rum runt en cirkulär reception.
Kvinna som spelar tennis i en ljus orange utstyrsel.
Fyra kvinnor stannar längs en gångväg för att titta på ett område bortom stängslet.
En indianfamilj som rider på en motorcykel på gatan.
En brun hund med orange krage hoppar för att fånga en färgglad boll.
Ett barn som leker med lite garn.
En parad av hejaklacksledare som bär svarta, rosa och vita uniformer.
En man i kostym hoppar mot sin brud.
Två officerare rider sina hästar längs en gata som gränsar till en grön och gul park.
En kvinna pratar med en liten flicka som spelar ett spel.
En person med rött hår och en svart skjorta står utanför, pratar och ger med händerna.
En person sitter på kanten av en klippa.
Två hundar tar tag i ett rött föremål på en gång.
En tennisspelare som rör sig för ett skott.
En man med tennisracket bär ett blått pannband och blå armband och spelar tennis.
En pojke träffar en tennisboll på en bana.
En tennisspelare springer på banan med sin racket i handen.
En pojke i en Mets jersey poserar på sin cykel.
Många människor sitter i en park och tittar på ett schackspel.
En hästkapplöpning på en gräsbana
Eleverna som sitter på gräset äter en lunch från en röd ryggsäck.
En pojke bromsar dansen som en publik tittar på.
Tennisspelaren gör sig redo att slå bollen som nästan är på honom.
En man i ett blått pannband som spelar tennis.
En person som håller i en tennisracket träffar en gul tennisboll.
Människor handlar runt ett utomhus system av butiker.
En liten pojke som bär en röd hjälm rider sin cykel längs en mönstrad stig.
Fotot är taget av två personer som går mellan bilar på en gata.
Ett par män som spelar gatuboll.
Fem personer har utsikt över den vackra staden.
Flera män i biofarliga dräkter bär en människoliknande docka på en rullande säng
En far släpper ut sin dotter i en pool vid Oceanside.
Flera unga pojkar spelar fotboll framför en stor brun trädörr
En grupp människor rider på sängen av en lastbil längs en grusväg.
En kvinna kramar en man vid ett kvällsevenemang.
Barn leker framför en stor dörr.
En vuxen man och en topless flicka dansar.
En flicka i rosa prickar tittar på en häst.
En flicka som bär hatt och håller en iPod sitter på sidan av en byggnad.
Två vuxna pratar medan ett moln av rök fyller bakgrunden.
Två personer tittar på en ljus utställning av något slag.
Gubben har glasögon, en halsduk och en hatt.
En pojke som utför ett väggtrick med sin cykel på en vägg täckt med graffiti.
En pojke har ett fiskenät.
En manlig tennisspelare som står på en tennisbana svänger sin tennisracket vid tennisbollen.
Två unga kvinnor, varav en är att föna håret.
En man klättrar upp för en sten medan andra väntar på sin tur.
Båtmannen jobbar på en ofullbordad båt.
En man använder ett verktyg på dessa långa träbitar.
Tennisspelaren spetsar tennisbollen på gränslinjen.
En klättrare med blå hatt är att skala en isig klippa.
Personen hoppar genom luften på skidor.
Två musiker, en kvinna i svart som spelar piano och en man i svart kostym som spelar flöjt.
Folk står och går på en loppmarknad.
En asiatisk kvinna är på ett marknadsstånd som säljer bananer.
En man gör ett stunt utanför på sin cykel
Ett barn i en röd och grå rock framför ett träskjul.
En brun och svart hund springer över det gröna gräset.
En liten pojke hoppar från en tegelvägg på ett bord nedanför.
Han sätter fötterna på ett skrivbord.
En man i blå skjorta bygger en båt ur trä i ett trångt arbetsutrymme.
En man som klättrar upp för istapparna på ett rockansikte.
En man i en grön tröja försöker skära något i ett kök.
En man som sitter på en veranda och säljer röda varor.
En kvinna som sitter på en trottoar med andra åt sidan och bakom henne.
En man med hjälm åker snöskoter.
Två hundar springer två en damm en vinterdag.
En brun hund som står i vatten.
Två cowboys repar en stut från hästryggen i en indoor corral.
En cowboy på en häst repar en stut.
Två små flickor på en studsmatta och en lekstuga är bakom dem.
Tre hundar leker i de grunda delarna bredvid en stenig strand.
Unga människor, både flickor och pojkar hoppar högt upp i luften på gatan de går ner.
Två personer går på en språngbräda.
Person med blå och svart kostym surfar.
En man och två kvinnor på en motorcykel.
En reparatör hänger ovanför en bredbilds-tv upphängd strax under taket i en katedral eller ett museum.
En man som står framför en disk och ser på en lagad mat.
En racerbil på ett spår har flammor som skjuter bakifrån.
Flera busiga barn leker med leksaksvapen i ett offentligt område.
En svart stor dansk som springer mot kameran på en bakgård
En man och en kvinna som sitter på stranden och tittar på landskapet
En grupp människor plockar upp något som brinner.
En hund ligger på ryggen på en väg.
En skateboardåkare rider en skateboard längs ett metallräcke framför en betongbyggnad.
En liten grupp människor sitter tillsammans utanför.
En grupp människor med en brandmotor i bakgrunden.
En kvinna sminkar en mans ansikte.
Två damer sitter i restaurangen och pratar och skrattar.
En judisk familj som har ett möte.
En tjej med vit skjorta och svart bälte dansar vilt med två kvinnliga vänner.
En grupp män går längs en väg delad med gula rep.
Fyra koreanska män sitter på en bänk och en av dem tar på sin mobiltelefon.
Hunden springer på ett fält.
En byggnadsarbetare som installerar ett fönster i en byggnad med en turkos dörr.
En man står och diskuterar med sina kollegor
En man sitter ensam och läser en tidning i ett fabriksrum.
Tre män med röda skyddsvästar står redo.
En man i hatt som håller i ett redskap står bredvid en häst som är fäst vid en släde fylld med hö i ett kuperat område.
En man som hoppar på väggen på en stor graffitivägg.
En grupp på sex personer sitter runt ett silverkonferensbord med anteckningsböcker och pennor.
Den här personen sitter på en tealbänk och läser en tidning.
En sjaskig hund springer nerför en grusstig i en frodig skog.
En man som håller i en gitarr och talar in i en mikrofon.
Konstnärer i vitt sträcker sig mot publiken.
En vitklädd man spelar gitarr.
Ett stort kryssningsfartyg passerar en strand där solbadare lutar sig under gula paraplyer.
Den grå hunden sitter tyst klädd i en blå banjacka.
En hund som försöker bita en man som tränar honom.
En kvinna som spelar softball har fångat en boll och faller ner.
En svart hund med blå krage sitter på beigematta.
En hund fångar en färgad boll medan han står i gräset.
Tre hundar racing på ett grässpår bär olika färgade tröjor.
En man som sover i en stol framför en full bokhylla
En flicka spelar en röd flöjt medan en annan tjej håller en rosa gitarr.
Två bmx ryttare racing på ett spår
Två kvinnor med mörkt hår står tillsammans utanför en buss.
Ett barn i en röd jacka som håller upp två fingrar.
En vit hund är pouncing på en brun hund i ett inhägnat i trädgården.
Två skäggiga män står bakom ett fall fyllt med cigarrer.
En stor lastbil parkerad nära ett garage som säger parfymer på framsidan.
Två hockeyspelare försöker få pucken.
Två hästar är fästa vid en vagn med hund och man inuti, och en kvinna står bredvid den.
Två kvinnor som rider i en motorcykel de båda bär hjälmar
Två personer i röda och vita uniformer på matchande randiga motorcyklar stannar i en plaza bredvid en hög vägg av betong trappsteg.
Tre män klättrar på varandra med gula och bruna skjortor.
En man i svart t-shirt hoppar något på sin orange cykel.
Flera människor väntar på sin tur att beställa mat.
En familj njuter av en måltid tillsammans, medan deras 4 hundar alla njuter av en tupplur på golvet runt bordet.
Två afrikanska kvinnor tillagar en måltid.
En brun hund som bär en rosa skjorta följs av en brun hund som bär en gul skjorta.
En vit pälshund springer genom löven.
Fyra män dansar på scen tillsammans.
Ett barn som håller en guldkanin stirrar på en P-formad kaka.
En basketspelare hoppar och ska dunka en boll framför en publik.
Ett barn i lila byxor springer.
En brun hund hoppar upp i luften
En svart hund som springer mot kameran.
En ung kvinna i grå skjorta sopar sin dörr med en kvast.
Mellersta Östern lagar mat i vita uniformer.
En gammal person sitter i en plyschstol med en stor vit hund som ligger ovanpå honom eller henne.
En liten hund springer med en brun boll i munnen.
Barnet bär en korg med färgade ägg och böjer sig över med ett ägg i handen.
Under ett basebollspel förklaras en Dodgers spelare vara säker.
Mat serveras till ett bord där en kvinna i en blå blazer sitter.
Två svarta hundar leker i snö.
En person som rider på en skateboard hoppar högt ovanför betongtrappan.
En grupp människor som står utanför en byggnad.
Kvinnan i blå outfit och stövlar står bakom lerig Toyota lastbil med ryggsäck nära buskar.
Cyklister håller sig i linje med varandra när varje person bär olika färgdräkter.
En brun hund hoppar över en röd ramp vid en agility park.
Två män med huvuden som skriver på en tidning.
En racerförare reser sig upp med handen pekande i luften.
Gitarriststrummor på scenen under strålkastarljuset
En asiatisk kvinna tittar på en svart jacka.
En äldre man köper mat på en asiatisk marknad.
Det finns ett äldre barn som rider en röd gummiboll fastbunden på ett blått rep och svingar från det.
En vandrare med ryggsäck vadar i en flod.
Ett ungt par sitter på en soffa och ler mot kameran.
Lille pojke njuter av en dag i parken
Två hundar, en ligger ner, leker på en gård.
En man som spelar fiol medan han läser sina musiknoter.
En kvinna sitter på en blå bänk framför en kullerstensmur mellan två träd.
Ett barn glider ner för en grön rutschkana.
En kille med glasögon och skägg i kostym är omgiven av fotografer.
Två pojkar tittar på en säl i ett akvarium.
En asiatisk kvinna i en röd lappad skjorta som bär två vattenmeloner nerför en trottoar.
Två personer fäktas.
En person åker skidor i snön, snön flyger bakom.
En man på en stenig topp.
Fyra musiker sitter i en halvcirkel på en scen och spelar sina stränginstrument.
Fem män i blå och svarta uniformer poserar för en bild.
En svartblå insekt som flyger över en vit blomma.
En äldre gentleman och en äldre dam pratar med två yngre damer i uniform på en stadsgata.
Gamlingen i hatt skär trä med en såg utanför.
En hund hoppar över ett stängsel.
En person sitter med ryggen mot en vit vägg med en brun hund.
En vit man som spelar ett instrument utanför.
En man jobbar med ett litet glassstånd som säger "Sorvette e Gelados" på sidan.
En matleverantör betjänar gärna sina hungriga kunder.
En man lutar sig åt sidan på en såpa racer mitt i ett hopp.
En ung asiatisk flicka sitter på marken i spillror.
En äldre kvinna läser en tidning på ett kontor.
Man gör kyssar ansikte för kameran, medan en annan man tittar på.
En flicka i rosa snödräkt stänker ner i smutsigt översvämningsvatten bredvid ett picknickbord.
Sju fotbollsspelare i en grön fält bär röda tröjor.
En kvinna skär av dreadlocks från en ung man med svart hår.
En man som sover på gräset under en grön filt.
Två personer rider en skidlift med berg bakom sig.
Folk går på gatan nära en jättelik tjurstaty.
En grupp människor står på en scen och håller färgglada hinkar.
En äldre kvinna som städar fönstret på en dörr.
Två män står på en klipptopp med utsikt över en sandstrand.
En kvinna i ett vitt förkläde balanserar en korg på huvudet.
Hunden springer med en gul boll i munnen.
Skateboarder i jeans och t-shirt som utför hopp.
Två män är inne och lagar mat över en eld.
Grupp av unga vuxna med hinkar och blöta våta på gatan.
En liten flicka i röd klänning och cape håller en stor tennis racket.
En man som tittar genom en kikare.
En person i grå snowboard nerför en kulle.
En man målar bredvid en byggnad.
En pojke i orange skjorta och blå jeans hoppar på rutschkanan medan andra tittar på honom
Tre personer sitter på en bänk under palmer.
Ett barn ler glatt när han håller fast vid en metallstång.
Pojkar på en fest som ritar på sin väns rygg med en svart markör.
Människor som äter vid ett långt bord fullt av mat och dryck.
Sex afrikanska barn sitter vid två bord.
Flickan har rosa byxor och en prickjacka på sig.
Folk går längs stranden en solig dag.
En pojke i en blå skjorta hammare på marken.
En äldre man står på kanten av en tågplattform.
En flicka i rosa kjol håller i en syster.
Två män sitter på en stollift.
En grupp människor har en stearinljus vaka till ära att rädda träd.
En gravid demonstranter håller upp en pro-Amerika tecken.
En man i jeans &amp; en cowboyhatt håller upp en skylt.
En man klipper en gräsmatta på en kommersiell egendom.
Muzzled greyhounds är racing längs en hund spår på natten.
En man i ryggsäck och hjälm som cyklar.
En mörk hund tävlar i en hundtävling.
Cykel racer nummer 661 vrak på smuts racetrack.
En pojke hjälper till att driva en ung flicka på gungan.
En ung flicka med grön t-shirt och blont hår.
En svart hund springer genom ett snötäckt område och håller något grönt i munnen.
Man åker snowboard nerför ett berg.
En man gör ett cykeltrick på en grusväg.
Två små barn leker gärna på en däcksvinge.
Två personer, klädda i långa dräkter, visas i en liten roddbåt i vattnet.
Mannen skateboardar över en stock i snön.
En man utan skjortskateboard på gatan
Unga vuxna som sitter i trappan och pratar.
En man som kör motorcykel när han bär svart uniform.
En man skär något ovanför ett handfat.
Flera människor runt en länsmässa med flera attraktioner inklusive en spådom maskin som kallas mormors förutsägelse.
En kille under vattnet i blå badbyxor som spelar död.
En byggnadsarbetare tar en paus medan han lutar sig mot en gul bar.
En ung man i brun jacka kör en rullande matvagn.
Ett litet barn i rött kastar en skiva.
Två smala vita hundar med två stående män i baseball kepsar
En stor, vit fågel åker skridskor över toppen av lite vatten.
En person i en röd jacka rider en mountainbike.
En svart hund i krage på andra sidan stranden.
Ett litet barn i grön skjorta är på en karusell.
Människor går förbi en ljus karusell; en del människor sitter.
En ung flicka som håller i ett uppstoppat grisleende.
Två flickor spelar på en uppsättning parallella barer.
En kvinna i svart och vitt är på cykel.
En kör i röda uniformer som sjunger framför ett företag.
En man och en hund leker med en gul boll.
En man med grå hatt som målar en scen av människor i parken.
Hunden flyr från kvinnan på stranden.
Brun hund hoppar över en bar på ett gräsfält.
En hund hoppar över en röd och vit grind.
En kvinna vinkar till folkmassan när hon rider berg-och dalbana.
En ung pojke sitter på golvet och sätter på sig sin sneaker.
En person som kör fyrhjuls ATV över ett hopp.
Ett barfota barn klättrar på djungelgymmet.
Ett barn som sover på betongen på någon sorts filt täckt med rockar.
En skateboardåkare i luften när du hoppar.
Brun och vit hund travar över jorden med träd i bakgrunden.
En motocross racer i grönt och en hjälm racing i smutsen.
En kvinna som håller i en mikrofon talar till en man i vit skjorta.
En skäggig collie hoppar över galler på en agility test kurs.
En man i svart hatt håller en liten flicka på sina axlar.
En ung pojke sitter i en grön tunnel
Den unga flickan svingar, och hennes hår flyger ut bakom henne.
En kille som åker nerför den snöiga sluttningen.
En ung flicka flyger en drake på ett fält bredvid många byggnader.
Man bowling i en svagt upplyst bowlinghall.
En ung flicka i skolan dansar uniform i en vattenskulptur mitt på ett trångt torg.
En ung pojke ramlar ner i en vattensamling.
En ung man sitter på en klippa och tittar på havet.
En barfota unge gör ett trick på sin skateboard.
Asiatisk baby som bär en tröja och sitter i en fåtölj och leker med en SvampBob leksak.
En rad åskådare på ett lopp.
Ett par människor rider ATV's på en grusspår.
Två män arbetar tillsammans med ett byggprojekt.
En man bär ett barn på axeln i regnet i en stor asiatisk stad.
En stad av by shoppare och åskådare njuta av den vackra dagen.
En kvinna i en vinröd kappa går ut Trader Joe's med en vagn full av matvaror.
Motocross ryttaren bär blå och svarta byxor.
En pojke knäböjer under en björnstaty som har en målning av en man på ryggen.
Tre äldre personer står framför en avrovulcan.com-skylt.
En kvinna som simmar i en pool blir plaskad av sin lagkamrat som simmar förbi.
En man klättrar utan utrustning.
Tre barn leker på en sväng i trädgården.
En flicka som flyter i havet en vacker dag.
En klättrare klättrar under ett överhäng högt över marken.
En cyklist hoppar på ramp täckt med graffiti.
En kvinna joggar medan hon lyssnar på sin iPod.
En pojke i blå kläder cyklar.
En pojke har vänt ryggen till i en simbassäng medan en annan pojke tittar.
En långdistansbild av en strand med människor och djur.
Två tjejer som leker klä upp sig och lägger upp den för kameran.
En ung man i en park förbereder sig för att fånga en frisbee.
En svart och vit hund leker i en damm eller bäck.
En kvinna ser en flicka leka i en stadsfontän.
Det är en ung man mitt i en komplicerad dans, och hans vänner hejar på honom.
En grupp människor poserar i ett konsertområde.
En man med glasögon och grå skjorta är på en fullsatt gata.
En cyklist i gul hjälm cyklar genom skogen på hösten.
Tre hundar springer längs en gräsbevuxen gård.
Tre vänner som hänger mitt i hoppet på en strand.
En flicka med vit ryggsäck står och mindre barn sitter i rad på marken.
En ung pojke ylar när en kvinna pratar med honom.
En folksamling samlas på ett torg.
Flera flerfärgade hundar springer genom gräset.
En man på en sele mitt i att klättra genom en grotta.
En kvinna håller ett barn i blått.
En pojke tittar genom luckan i ett rött och vitt tält.
Man med fjäderfä på ett bord.
Män i kamouflage byxor racing över en parkeringsplats.
En rödhårig flicka hoppar av en svan.
En man i svart väst och vit knapp-up sitter med en kvinna i en randig tröja.
En hund springer under en tävling.
En ung blondhårig tjej får sin frisyr av någon i en gul blus som håller en vit kam.
En man hoppar över en brun stol medan han skateboardar.
Racing bil märkt TEAM PENSKE på spår, banderoller och åskådare i bakgrunden.
Folket har färg på sig.
En kvinna i orange skjorta tittar upp på en man som står på en balkong.
En man och kvinnor som sitter på en restaurang eller bar.
En hukande vit man i gul skjorta ser ner från toppen av en trästruktur.
En lärare som hjälper en elev på en datorstation.
En man i shorts går en stor brun hund och en kvinna som knuffar en barnvagn går precis bakom honom.
Två barn i en flotte på en vattenrutschbana.
Ett barn i lila kläder leker med en leksak inuti en gård med andra leksaker och ett staket.
En kvinna går en barnvagn på en pittoresk stig.
Det finns 2 män klädda i ränder som sitter under ett grönt paraply.
En kvinna fotograferas när hon står bredvid ett konstnärligt monument.
En brun hund som springer på stranden nära havet.
Den här personen städar byggnaden med en grön hink.
En man låter en tandläkare undersöka tänderna.
En kvinna sitter på en sten vid kanten av ett vatten.
En nobbad hund i ett lopp, med fyra hundar efter.
Tre män sitter på golvet i grönt rum.
En publik ser en grupp elddansare uppträda.
En man som hoppar ut ur en helikopter i havet.
En grupp pojkar sitter nära trottoaren och två ler medan en gör ett ansikte.
En brun hund galopperar genom gräset.
Barn som tittat igenom tidskrifter de har vika in i rör
rugbyspelarna spelar på en plan.
En ny brud klädd i vitt kastar en bukett till väntande kvinnor bakom henne.
En tävlingsbil med ett moln av damm bakom sig
Två vuxna ställer sig på en buss och tittar ut genom fönstret.
En man i brun jacka står på en buss.
En grupp artister sjunger och arbetar för att underhålla publiken.
Två män med solbrända hattar som arbetar i en trädgård.
En man i blå jeans, vit skjorta som drar upp en lina ur vattnet.
En blond kvinna på stranden som hoppar runt när hon njuter av sin ungdom och frihet.
En skara människor är vända åt samma håll medan somliga håller sina händer i luften.
En båge gör ett trick på sin skateboard i en skatepark.
Det här är en liten flicka som står framför en glidbräda och blåser bubblor.
En pojke som bär hörlurar poserar i köksdisplayen
En man i röd skjorta, med två kvinnor och en annan man som står på någon sorts marknadsplats.
En man hugger en tjur i en tjurfäktning.
En man som gör ett trick i luften på sin cykel.
Lilla flicka med stickad mössa, doftande blommor.
En man i skjorta sitter på lekplatsutrustning.
Folk stannar för att ta in landskapet på bron.
En man står på passagerarsidan av en svart bil.
Två hundar tävlar över ett fält en solig dag.
Flickan klädd i rosa och vitt, och bär en stickad mössa, sträcker sig mot ett blommande träd.
Folk sitter runt ett bord med mat.
En kanna på en kulle kastar en baseball.
En liten flicka leker nära en höbal.
En liten flicka i grå skjorta ler när hon borstar tänderna med en gul och orange tandborste.
En svart och vit hund som springer från under ett gult täcke med en person bakom sig.
En grupp människor i blå kläder slappnar av på gula maskiner.
En man står bredvid ett gult fordon.
Denna familj behöver vila efter sin långa promenad så de stannar vid parken för att mata duvorna.
En kvinna och flera män bär ansiktsmasker på en tunnelbana.
Två män brottas på en blå matta.
En tjej i grönt hoppar på betong.
Tre basebollspelare i rörelse; en glider in i en bas, en annan kör i bakgrunden.
Här är unga pojkar som åker skridskor på en tjänsteresa.
Ett litet barn i vit och gul utstyrsel sträcker sig efter ett gult papper japansk lykta på ett trästaket.
En hund som springer på en strand.
En liten flicka med en gul klänning som gungar i en liten vit stol.
En kyrkosammankomst lyssnar på en körföreställning.
En person i gult är att cykla på en grusväg.
En brun hund bär en lång käpp på det gröna gräset.
Tjejen med blå skjorta springer genom ett vetenskapscenter.
En kvinna som sitter på en bänk och läser en bok.
Sju flickor utgör en gruppbild, med tre flickor som bär slips, och fem flickor som bär klänningar
Arbetare på Basking Robbins är väldigt upptagna.
Ett gäng killar i svart spela paintball.
Landhockeyspelaren tar en grävare i en match.
En kvinna som bär en orange väska går nerför gatan med sin vita hund.
En man och en kvinna joggar längs trottoaren.
En asiatisk kvinna håller upp sina händer och flickan bredvid sina klockor.
Två män sitter bakom en glänsande svart disk med matchande svarta kostymer och lila skjortor.
En grupp människor står runt dj utrustning inklusive en skivspelare och en ljudmaskin.
En kvinna i en ljusfärgad klänning sjunger för en publik.
En tennisspelare i vit skjorta slår bollen.
Mannen i shorts serverar tennisbollen.
En kvinna med vit t-shirt och svarta shorts är på väg att träffa en volleyboll.
En kvinna bär en volleyboll.
En man i solglasögon och en basebollmössa hoppar för en gult randig volleyboll.
En man på en mountainbike utomhus.
En man som bär skjorta och slips, ser förbryllad ut när han navigerar genom en folkmassa.
En svart och brun hund som tittar på en fluga.
En man och kvinna pratar på en utomhus loppmarknad där konst visas upp.
En tjej med pannband bär en rosa skylt på gatan.
En man med en ovanlig frisyr i en t-shirt bär två tallrikar mat.
En man med grön skjorta och vita shorts spelar volleyboll.
Många människor samlas och gruppen i förgrunden samtalar med drycker och deras kylare i närheten.
En snowboardåkare gör ett trick på en halv pipa.
En man cyklar genom gräs i ett skogsområde.
En man mountainbike med blå hjälm
En man i gul utstyrsel tävlar sin cykel i vildmarken.
En grupp människor står och väntar på att få se något.
En man tar en bild av ytterligare två män i en folksamling.
En kvinna i grå skjorta sträcker sig i en utomhus parkområde.
Arbetare i västar och hårda hattar arbetar på gatan i en livlig stad.
Tre män står i ett glasområde.
Ett barn som är klädd i blå skjorta och mössa bär en fotbollsboll.
En liten flicka i en hatt som klättrar på en barnvägg.
En man med glasögon hs mat i händerna.
En man som målar en stadsscen.
En flicka står på gräset och håller i en rullande låda med en vit hatt på gräsmattan och solglasögon.
En man i brun skjorta, hade och axelväska stående med två kylare.
En man och kvinna är i köket och ett paket Challengesmör ligger i förgrunden.
Människor i hemgjorda kläder sitter vid skrivbord.
Tre små barn och en kvinna paddlar nerför en flod omgiven av tjock vegetation.
Ett band uppträder på scenen.
Fotbollsspelare samlades alla på ett fält för ett spel.
Den stora svarta hunden är bakom den lilla svarta hunden.
En pojke som bär en röd skjorta på en skateboard hoppar upp för några trappor
En bicyklist utför ett trick på ett högt träd.
En grupp barn leker på en däcksväng.
En grupp människor vilar på en järnväg i ett köpcentrum.
En försäljare, som bär en storbröstad solhatt, sitter på en pall bredvid sina varor.
Flera människor sitter och slappnar av i snön.
En skateboardåkare fångar stor luft vid skateparken.
Den lilla flickan bär rosa är att ha kul bungee hoppning.
Den svarta och bruna hunden rullar i gräset.
En kinesisk restauranganställd som ger en matverkstad.
En ung kvinna som läser ett nummer av tidskriften People.
En kvinna hoppar med armar och ben utspridda nära en bostad.
Två män fiskar flugfiske i en låg murkig damm.
Två unga pojkar brottas medan en vuxen man tittar på.
Två flickor dansar och en har papper i handen.
En svart kvinna som jobbar på en fiskmarknad.
Det här bröllopsfotot visar bröllopsfesten, i lila och vitt, som samlats utomhus.
Två hundar tävlar på ett spår.
Pojken bär blå solglasögon och hoppar förbi en gul räcke.
En man jagar en motståndare i en rugbymatch.
En dansare på en scen utför ett drag som involverar hennes meddansare som står bakom henne och sticker ut sina armar så att det ser ut som om hon har flera armar.
En kvinna spelar ett musikspel i en arkad.
En kvinna med solglasögon på huvudet och stående framför en konstutställning.
En äldre man sitter vid sitt skrivbord, som står framför en butik och läser kort.
Två barn leker på ett fält av röda blommor.
Tre välklädda barn sitter på en bänk och ler.
En man som drog två barn på en släde på en snötäckt väg.
En rodeo ryttare rider en häst på en arena.
En flicka i rosa kläder tittar igenom bagaget i en tältstad.
En man som navigerar en vattenfarkost under delvis molnig himmel.
En äldre kvinna går förbi en vägg med hjälp av en käpp.
En grupp flyktingar som sitter bredvid sina tält.
Två soldater går in i ett tält med män och kvinnor som bevakar dem.
En svart pitbullhund springer genom jorden.
En man går på en slingrande gata med en regnbåge i himlen.
Två motorcyklist racing runt ett spår
En clown med färgglada byxor som sitter på en bänk i en gammal byggnad.
En surfare fångar en bra stor våg.
En man är nära vatten i en stad och är klädd i våtdräkt, snorkelmask och hjälm.
En man som tittar åt vänster och går nerför gatan.
En pojke rider en scooter ner för betongvägen.
En grupp barn håller i ett rep.
Två män hoppar från ett picknickbord, med en klippvägg och skog i bakgrunden.
En ung flicka som blåser på en maskros.
En liten flicka i blå skjorta går ensam på en gul parkeringsplats.
Folk håller pappramar framför sina ansikten.
Fyra tjejer dansar i matchande kläder på en gatufestival.
Två hundar springer över den karga marken.
En person i en vit hjälm står bredvid en stege.
Vissa människor är klädda i klassisk europeisk klädsel, medan de håller böcker och en trumma.
En asiatisk man med svart hatt håller en liten asiatisk flicka i sina armar.
En hund ligger på rygg med en favorit tennisboll i munnen.
Spelare i röda uniformer på bänken under en hockeymatch.
En kvinna hoppar över ett hinder under ett lopp.
Ett naket barn kryper på stranden framför en häst och en man.
Två små barn med långa ärmar står i gräset.
En liten hund med en leksak i munnen hoppar över en påle.
Två män under en fotbollsmatch
En ung flicka leker i en källa med vatten.
En tjej som spelar softball slår till.
Den första baseman dykning för att fånga ett kast, medan löparen berör första basen i en softball spel
Tre personer spelar baseball på ett fält i en park.
En kvinna och två unga män som står varandra nära.
En flicka kliver av kullen efter att ha kastat den första planen ut på en basebollmatch.
En kvinna som äter med ätpinnar sitter framför slaktat rått kött.
En man som tittar ut på baksidan av sin bil och tittar på en gul skåpbil bakom
En koppelhund är på bakgården till någons hem.
Två svarta hundar leker i gräset.
En rugbyspelare i svart trycker sig igenom en spelare i rött medan han bär bollen.
Tre män som bär rutiga skjortor skär trä.
En restaurangarbetare med orange skjorta som sätter ketchup och senap på smörgåsbröd.
En snowboardåkare som gör ett enhands armstöd.
Tre barn sitter högst upp på en trappa.
En blå Subaru rally bil vänder ett hörn med åskådare.
En brun hund och en svart hund som slåss på en inhägnad gård.
En man och en pojke leker i sanden.
En man i läderrock tittar in i restaurangen och tittar på 2 tjejer.
En brun hund på gräset bredvid en damm.
Två vuxna par satsar på ett kasinobord.
En kvinna i gröna skridskor genom en gatumässa.
Ett litet barn toppar huvudet bakifrån ett stort brunt paket.
Folk tittar på en racerbils hastighet.
En mörkbrun hund hoppar bakom en ung flicka i shorts.
Äldre kvinna med klyvning sätter på mascara förföriskt i spegeln.
En ensam cyklist som hoppar på sin cykel framför en graffitivägg.
En delfin sticker över vattnet.
En ung dam gör ett köp från en man med en push cart.
Man i randig skjorta med handskar på svetsmaskiner.
Fyra personer i ett växtfält, bakgrunden verkar vara i Indien.
En man dricker apelsinjuice och går ut.
Ung blondhårig, blåögd pojke spelar på en repbana på en lekplats.
En liten unge med en gul och röd fotbollsleksak.
En grupp arbetare är på ett åkerfält och planterar vete för året.
Ett band bestående av en kvinnlig basist, en manlig ansiktsmålad gitarrist, och en medelmåttig sångare på scen.
En man som håller ett barn och ler, sitter i bänkarna i en kyrka.
En kanna som bär nummer åtta går igenom pitching-rörelsen.
En umpire tittar noga när en vänsterhänt kastare kastar en pitch från högen.
En ung kvinna med en rosa mask över ansiktet.
Ett barn i gult och svart sparkar en blå och svart boll.
Några afrikaner som leker med en boll.
Två racerbilar kör fort på ett spår med rök som kommer från baksidan av dem.
Två hundar på stranden, sprang i vattnet
Fyra män leker på ett stenlagt område.
En äldre man sparkar ett föremål.
En brun och vit hund framför ett skjul överväldigad av angrepp av tennisbollar.
En man är på ett litet drag längs trailer arbetar med landskapsarkitektur material.
En figur av en orientalisk man sitter på en vägg framför några vita hyreshus.
Tjej med svart färg under ögonen går, flicka i förgrunden av foto.
Hon målar en gul blomma på vitt papper och övar på att bli konstnär
Äntligen fick han en bar på sin wifi-anslutning.
Två män sitter i rundade gröna stolar på ljusblå matta.
En kvinna som beskär en prydnadsbuske på sin gård.
En man har en trofé på scenen.
En man äter utomhus med en grupp människor.
Tre kvinnor och två män i baddräkter, sola på gräsmatta stolar täckta av handdukar.
En man använder en kvarn på ett skåps lås
Två mindre hundar jagar en större hund runt en damm.
Pojke i gul skjorta får bilden tagen omgiven av duvor
Tidsfördröjning foto av två barn som leker i en pool av vatten.
En ung flicka som håller en docka ler.
En man och en kvinna står knäna djupt i de hårda vågorna bredvid en röd-orange båt.
En man kör en röd racing motorcykel.
En manlig surfare i luften, lämnar vattnet.
En pojke som sitter på golvet och tittar upp på en kvinna i en grön stol.
Tre personer och en hund står framför en flod en kall dag.
Två kvinnor spelar tennis.
Två sjukvårdspersonal tar hand om en patient och tar hänsyn till hans eller hennes journal.
Den unge mannen sparkar en fotboll på dammig mark.
Tre män i en klar orange båt ras över vattnet som skum sprayer i luften.
Två hundar leker boll tillsammans utanför.
Två personer flyttar slangen när andra arbetar i trädgården.
En grupp människor går nära några träd.
En man i våtdräkt på en surfbräda.
En grupp människor låg i skuggan.
En grupp tjejer med en i blå skjorta med ryggen mot kameran skrattar.
En man som står på ena foten med en liten flicka framför en katedral.
En ung man ställer sig i kö i footballträningen.
En fotbollstränare och fotbollsspelare som tränar.
En man sitter på gräset och försöker få ett hål i en fisk.
En kvinna i lila leggings går tvärs över en gata.
En man som ser ledsen ut med renare och ett verktyg bredvid sig.
En brun labradoodle hämtar en tennisboll i en sjö
En asiatisk man navigerar en båt med 2 passagerare nerför vad som verkar vara en flod djupt inne i skogen.
Ett par cyklar för två.
Den lille pojken har jätteroligt i vattenparken.
Två män och ett barn som arbetar utomhus med olika utrustning.
Man i vit skjorta och bruna shorts gör ett trick på en skateboard.
En ung pojke läser en tidningsbok utanför.
Ett barn hoppar på en uppblåsbar dörrvakt.
Surfaren rider en våg med ett berg i bakgrunden.
En komplex byggnad ligger i bakgrunden med människor som står runt och några cyklar.
En kvinna som skriver medan hon står vid männens sida.
Många asiatiska kvinnor går ut i ljusblå skjortor.
Flera män runt en inomhus basketkorg.
Man i ärmlös skjorta och shorts står i mitten av golvet.
En man hoppar in i en mörk gymnastiksal.
En grupp män står i en gymnastiksal med en basketboll.
Kvinnan poserar i höga klackar på en rostig stege.
Asiatisk man klädd i vitt, med halmhatt och handskar, som ger sig på folk i mängden.
Två gatumusiker spelar gitarr i Asien.
En man med vit och röd hatt spelar golf och kommer att försöka träffa bollen.
En grupp människor poserar med sina hundar.
En grupp människor går på gräs nära en sjö med hundar som leker runt dem.
Två unga kvinnor med ett stort papper.
Många löpare springer på gatan i ett lopp.
En gulskjortad löpare springer med ett nummer fastsatt på skjortan.
En kvinna med svart skjorta tittar på en karnevaltur.
En man går förbi en latinamerikanska fabrik.
En stor grupp människor går på en trottoar.
Hund simmar genom vatten bär käpp i munnen
En pojke slipar ner ledstången på en trappa med skateboarden.
En grupp människor bär siffror på gatan.
En rugbymatch pågår visas med domaren tittar.
En pojke som cyklar medan en man håller i cykeln.
Två oxar som springer genom sjön lämnar människan bakom sig, täckt av lera.
Fyra personer använder musikinstrumenten.
En hona hjälper ett barn att köra en stötfångare bil.
Människor som står runt ett torg med cyklar.
En man går nerför en gata av en man som säljer saker ur ett bås.
En surfare rider en våg när den kraschar på stranden.
Ett par sitter på en lutande trädstam och poserar för kameran.
En fotbollsspelare är att tackla spelaren med fotboll som publiken klockor.
En överbefolkad buss som reser nerför gatan med folk hängande på baksidan av den.
Tre personer som håller sig borta från solen
En grupp barn som sitter på golvet i ett konstmuseum och lyssnar på en äldre dam.
En svart hund som leker med en lila leksak.
En grupp rullskridskor på en sluttande väg.
Två motorcyklister tävlar runt ett cirkulärt spår.
En ung flicka spelar "kike-a-boo", som täcker ögonen på mannen på vars axlar hon sitter.
Sju personer hoppar ner i vattnet.
En kvinna som bär en T-shirt och shorts går förbi en röd Sedan
En man i blå mössa arbetar med en rosett.
En kvinna i vit skjorta och jeans som håller två krattor när hon går nerför gatan.
Rollerblader i röd skjorta åker skridskor på en ledstång.
En asiatisk temarestaurang med stor monterad fisk.
En man lutar sig mot en racing motorcykel.
En äldre man använder sin käpp för att peta i ett hål i marken.
Två kvinnor sitter på en parkbänk och pratar med varandra.
Ett barn i grå rock som sparkar en fotboll.
En brun hund hoppar över ett stängsel.
En grupp på cirka 11 personer i alla åldrar med kikare i skogen
Pojkar och flickor i marinblå skjortor ler för kameran.
En kvinna ser en hund hoppa nerför trappan.
Ett barn i Musse Mouse-skjorta har armarna uppe och verkar hoppa.
Ett barn i en blå jacka tittar till vänster när cykeln rider nerför gatan.
Skidåkaren åker nerför ett stort berg.
En kvinna klättrar uppför ett brant berg över vatten.
En man avfyrar ett vapen på skjutbanan.
De två hundarna står med huvudet sammanflätat runt varandra.
En grupp åkare är på en skatepark.
En man i skyddsväst som cyklar på motorvägen.
En man går på en fin trottoar bredvid en övergiven bar.
En manlig bicyklist som försöker få något från sin ryggsäck på en livlig gata.
Pojken hoppar sin cykel upp i luften.
En asiatisk kvinna cyklar medan hon bär en respiratormask.
Damen bär en bandanna runt hennes ansikte för att skydda henne från damm.
En kvinna med röd hatt och ansiktsfärg ler mot en annan kvinna.
Barnet leker i klippan.
En kvinna i en brun topp med glasögon står framför ett diagram.
Tre unga svarta män lutar sig tillbaka mot en vit jeep.
En grupp cykelförare som bär hjälm stående nära en skåpbil.
En trumpetspelare spelar musik med sin partner.
Två kvinnor tittar på en matförsäljare, med tanke på om de vill köpa något.
Ett litet barn som klättrar upp för stegen efter någon.
Polisen i ljusgula jackor tittar på publiken.
En man använder sin dator i ett kök.
En kvinna som bär en röd och vit klänning håller händerna med mannen i en blå jacka med blommor på sitt knä.
Flera män laddar en metallkanon
En kvinna i brun skjorta pratar med någon.
En kvinna presenterar olika dokument med hjälp av multimediautrustning.
En ung flicka är på en åktur på en nöjespark.
Två män står framför en stor grön lastbil.
En familj går genom ett grusfält under högbyggda träkonstruktioner.
Två svarta hundar tävlar om en boll på stranden.
En kvinna i en blå topp jobbar på en fabrik.
Fotgängare och en cyklist rör sig lätt förbi en modern byggnad.
Två tjejer leker i duschen med kläderna på.
En kvinna håller ett barn i armen medan hon pekar.
Det är en svart hund som hoppar in i en simbassäng.
En man kör en gruscykel över en kulle.
En man står mitt ibland en skara människor medan han röker en cigarett.
Fem män som släpar i ett fiskenät på stranden.
I en tom, dimmig bowlinghall förbereder sig en kvinna för att släppa en röd bowlingboll mot en grupp på fem stift.
En flicka som bär rosa svänger över en bäck.
En dam med lockigt brunt hår står i en publik med en kamera.
Två unga fotbollsspelare tävlar mot målet.
En grupp små barn i rullstol drar varandra genom en liten by när de fotograferas.
Äldre man leder bandet när de spelar.
En man i rutig gul med två tennhinkar.
En man som går en stor svart häst.
En smutscyklist tar ett stort hopp i gul kostym.
En hemlös man går ensam på trottoaren.
Ung pojke med en Elmo t-shirt som knäböjer vid ett bord med sin måltid.
En liten pojke ligger i en hög löv bredvid en skateboard.
Två softball spelare försöker fånga en boll
En dam kör sin hund genom en smidig kurs.
En bit kött presenteras ut genom fönstret i en butik medan en ung man går mot den.
En man som rakar sig med rakkniv.
En folkmassa står framför en byggnad medan de håller tidningar och håller flaggor.
Tre tjejer med huvudomslag som bär föremål medan de står på obelagd yta.
Ett par sitter på en parkbänk med lila ballonger bundna till den.
En tävlande i hästryggssvärdsstrider. Publiken ser på.
En kvinna som bär handväska går förbi en affär.
Två hundar springer på ett fält.
En dam som står vid disken på ett bageri och ler mot kameran.
Farfar, far och två söner sätter ihop ett pussel.
En grupp män i vita hattar inne i en industribyggnad med en som fotograferar en bild.
Män som står på en byggarbetsplats.
Den svarta hunden drar i något lila med munnen.
En liten pojke som bär en liten flicka på ryggen.
Fem personer står på en scen, gör sig redo att uppträda, som är oigenkännliga på grund av bristen på belysning.
Många individer med täcken på huvudet trängde sig samman.
En grupp män omger en kvinna i en slöja.
En ung flicka som står ensam i en hall.
Den söta lilla flickan med den röda borsten kammar håret.
Två arbetare i orange västar går med lastbil och riskkottar.
En flicka och en kvinna poserar medan de sitter i en mattad trappa.
En spelare glider in i hemplattan med catcher vakta den.
Två kockar, en i traditionella köksdukar, den andra i kostym lagar asiatisk mat i woks.
En smet gungar på en boll.
En högtidlig ung man i en randig krageskjorta håller en bild av sig själv och en kvinna i en silverram.
Chef med två kvinnor som har ett samtal.
Svart och brun hund hoppar över hinder med vita stöd.
Kvinnor och små flickor som utför en kulturell dans.
Unga flickor uppträder ett dansnummer på scenen.
En grupp pojkar som studerar i ett bibliotek.
Två unga asiatiska flickor klädda i något slags gröna och gula kläder dansar tillsammans.
En basebollspelare fångar bollen medan smeten når basen.
En kvinna med långt hår fångar en softball i ett softballfält.
Lilla flicka och äldre man, håller hand och går på tågspår.
En kvinna som håller en handdocka framför en klass av elever.
En hund hoppar för att fånga en boll i surfandet.
Två män klädda i gula uniformer använder en jackhammer i marken.
Två män i badbyxor står på sand.
En hund som jagar en tennisboll över ett gräsområde.
En äldre man som hänger sig åt en flaska bärnstensvätska.
En mamma knuffar sina två barn på gungan.
En man utför en smuts cykel stunt över sanden.
Spelare som bär orange, vit och svart jackor och några av dem pratar med varandra
En hund med en orange boll i munnen som simmar.
En pojke lutar sig ner framför en flicka med blått randigt hår på en tunnelbanestation.
Någon surfar under en våg på en vit surfbräda.
En softball spelare i rött och vitt gungar och träffar den gula bollen.
En flicka i röd och vit uniform svingar ett slagträ.
Två spelare är på ett vått fält och en är på marken.
En grupp tonåringar samlas på balen.
En ung pojke på en skateboard gråter medan en vuxen rör vid hans axel.
Hon är på väg att kasta en pinne för en tävling.
En tjej med rörigt hår har huvudet på pojken som ligger bredvid henne.
En person som hoppar en häst över ett stängsel.
Kvinnan hoppar en lång sträcka medan folk tittar.
Man rider på cykel när andra går.
En liten flicka i lila tröja och enkla shorts går med en kvinna förbi en tunnelbana.
Föräldrar tittar på när flickor spelar softball i ett spel.
En tjej som bär nummer ett LaFayette softball uniform är på väg att kasta bollen.
En tjej i vit och brun uniform svänger på en softball.
En softball spelares lag tittar på när hon svänger på en pitch.
En ung flicka förvränger sin kropp under en föreställning.
En ung flicka blåser bubblor med en orange bubbla trollspö.
Två killar som skojade med varandra.
En man står på en mobiltelefon framför en filmaffisch.
Tonåringar som bär formella kläder står i en grupp utanför.
En kvinna i blått står med en hand på en torr stenyta.
En skateboardåkare går nerför några trappor.
Två män går nerför en stentrappa, en åker enhjuling.
Många människor går genom ett shoppingområde på landsbygden.
Ett litet barn klädd i grön rock, blå jeans och rosa stövlar kastar sand på havet.
En person som tar en bild av en grupp andra människor.
En kvinna klappar sin hund nära en stenväg.
Den bruna hunden springer på gräset.
En man som står framför två annonser förbereder sig för att kasta något över ett fält.
En liten katt som ligger med en stor hund
Tre personer står framför en blå vägg med graffiti på, medan tre metallstolpar och tre gröna lådor är i förgrunden.
Hund med öppen mun och en leksak i närheten i luften
En grupp människor sitter i en hörsal och tittar på en skärm på scenen.
En man med svart hatt och glasögon som spelar gitarr.
En pojke i röd skjorta tittar mot en staffli som en konstnär har.
En man i supermankostym håller ett tecken på vägen.
En man och en hona lagar snabbt till ett däckrör på jorden.
En pojke som hoppar från en gul vårbräda.
En gyllene hund tittar på en blå och gul leksak på gräset.
En manlig artist spelar cello.
En ung, välklädd svart man som satt bakom ett trumset och log.
En kvinna med glasögon tittar på mat.
Två tonårsflickor sitter vid ett träbord och skapar hemgjorda hantverk.
En kvinna som kliver ur en röd flygande bil.
En blond kvinna vid ett bord skriver i en bok när två män tittar på.
Mannen i svart skjorta gör sig redo att kasta bollen i bowling gränd.
En flintskallig man i en blå blazer i en bok vid ett skrivbord framför en kritbräda.
En kvinna och en ung pojke.
En man i blå skjorta går framför en affär på en gata.
Två militärer utövar en "nedtagnings"-manöver.
En liten flicka hoppar upp i luften bredvid en jukeboxmålning.
Några går nerför gatan.
Två personer sitter på en träbänk och möter varandra för att prata.
Fyra vuxna som sitter vid ett bord och äter en måltid
Fem stora hundar springer genom en inhägnad gräsyta medan de bär mynningar.
Två små barn slår på en bongotrumma.
Surfare delvis synlig genom kraschande våg, stranden i bakgrunden.
Crowd tittar på flygplan och helikopter i himlen.
Ett barn cyklar högt i luften.
Ett barn som klappar en hund.
En grupp pensionärer sitter vid runda vita bord medan de väntar på mat.
Spelaren sparkar en fotboll på gräsfältet.
En grå hund och en solbränd hund som leker på ett gräsfält.
Sju sjömän klädda i blått på en båt.
En kvinna tittar genom ett vetenskapligt instrument på en liten bit teknik.
En man i en blå t-shirt håller en kamera.
Gruppen av människor gör enstaka fillinjer på fältet.
En man som sitter i en blå metallstol.
En hund med en käpp i munnen som går genom vatten.
En elev klipper papper med glädje.
En svart hund i en bandanna springer längs en grusväg.
Hockeyspelare rör sig snabbt mot pucken.
Skateboarden faller ifrån skateboardåkaren när han försöker hoppa.
En brun hund som leker med bubblor.
Två män i svarta uniformer som pratar med en man som håller i en flaska läsk.
En del män och kvinnor dricker vin medan de tittar på TV.
Period re-instruktörer sitter på gräsbalar och pratar medan andra i modernare klädsel sitter och går i bakgrunden.
En kvinna i en rutig skjorta som tittar i en glastank.
Folk sitter, står och läser tidningar i en gränd.
Baseballspelare med slagträ.
En kvinna i gul jacka och brun hatt står på en stig vid en sjö.
Vandrare går längs en tuff terräng.
En man med spade gräver i ett hål utanför.
Två äldre män i rockar står utanför.
Den lilla bruna hunden springer förbi en annan hund på gräset.
En fågel flyger lågt och vingarna breder ut sig.
Folk ser på när en kille tar hand om en fast växelcykel under ett tält.
En stor park bredvid en vattenförekomst med stora djurskulpterade buskar.
Två leende flickor står på en grusväg i Indien.
En brunhårig flicka går och hämtar en liten vit valp på en tom gata.
En blond kvinna i röd kostym som städar ett metallföremål.
Fyra hundar springer på ett fält.
Tre personer som håller i kameror står på en grusstig med gräs på sidan av den.
Äldre kvinna i orange klänning står på en strandpromenad.
En fet man i lila skjorta som äter ett potatischips.
En kvinna i rosa skjorta undersöker sin kamera.
En man vid namn Luke, som bär en ljusblå skjorta och en namnskylt, fotograferas från toppen medan han står lutad mot baren.
En man med en hund står utanför på tegelstenar och håller ett tecken.
En kvinna använder en symaskin på ett rörigt bord.
En äldre man går förbi och skriver på en vägg.
En liten svart och vit hund som bär en röd hink i munnen
En man med hjälm står framför en byggnad
En hane gör ett öppet ben trick medan han gör en wheelie på sin cykel.
En kämpe ger ett hårt slag mot ansiktet på en annan kämpe.
Två manliga UFC-kämpar boxas mot varandra i en ring.
Flera människor rider kamel 2 per kamel i öknen.
En kvinna i rosa njuter av sitt iste och aptitretare på en restaurang.
En skara människor som setts ovanifrån, flera håller kameror.
En kvinna och ett barn som försöker spreja en cykel.
En pojke på en cykel hoppar över några sandhögar.
En fotbollsspelare är på väg att fånga en fotboll.
En grupp människor sitter runt ett skrivbord.
En tjej som försöker träffa en boll i luften med en tennisracket på tennisbanan.
En pojkskateboard på en ramp.
En fantastisk outDoors Cafe på en solig dag.
En kvinna tittar på ett fotografi.
En man i hjälm gör stunts på en cykel.
Joggare springer längs en landsväg i ett lopp.
En brun hund dricker vatten från en skål medan en svart hund hoppar ner bredvid honom.
En hockeyspelare bär en röd uniform sträcker sig för pucken som andra följer.
En man sitter i en stol och tittar på en lavalampa och en datorskärm.
Två cyklister, en med mask, poserar på gatan med sina cyklar.
En skidåkare som hjälper en skidåkare att komma upp från snön
Pojken i röd och vit kostym är på en skateboard.
En man som cyklar nerför en ramp mot en smutscykelbana.
Mannen i skelett-tryckt läder outfit sitter astrid en röd motorcykel.
Två män pratar med en annan man som bär en blå mössa och bär en bok.
Ett par övar olika sätt att bära solglasögon framför en röd bil.
Män cyklar samtidigt som de försöker bära föremål framför en blå byggnad med röd trim.
En showgirl sätter på sitt läppstift i spegeln.
En bmx mc är för närvarande i luften gör en front flip.
Hockeyspelare som spelar hockey under en match.
Hundar tycker om att jaga varandra i parken.
En man med grå skjorta med vit namnbricka.
En man står mitt emot en kvinna och håller sitt halsband medan hon tittar på honom.
En liten pojke är i ett däck
Folkmassorna står runt omkring några palmer på jämna timmar av natten.
En leende man på en häst framför borste och skog.
En man och ett barn står på en gård bredvid en bänk.
En liten pojke gör ett handstånd på ena handen.
Ett rum fullt av barn lyfter händerna, fingrarna utsträckta, mot himlen.
En ung flicka poserar med en annan kvinna varje leende.
Tre unga vuxna tittar på den annalkande stormen.
Tre barn sätter sig ner till en måltid.
En man hoppar högt och håller flera blå ballonger på ett snöre.
En grupp barn sträcker sig på färgade mattor.
En man och en kvinna är fastspända i en rund metalltur.
En rugbyspelare blockerar medan han håller bollen.
En man i silverrock och hatt sitter på en buss.
Två flickor ger fredstecken.
En man står bredvid en kvinna och håller en elektronisk apparat i örat.
Tre seniorer tittar ut genom fönstret vid vattnet.
Folk passerar genom staden medan en musiker spelar.
Två personer står utanför en röd bil i staden och kramas.
Två kvinnor går nerför trottoaren vid en damm.
En kille som dukar bordet till middag.
En liten flicka i rosa klänning som håller i en slang.
Två hundar närmar sig varandra i gräset.
Ett antal människor sitter på en restaurang medan en servitör navigerar mellan borden.
Barn leker runt lekplatsen fartyget med klätternät och trappor.
En vit man, en svart man med röd halsduk och en blond kvinna som röker.
Gamlingen spelar dragspel i ett gathörn.
Elever i ett klassrum av något slag gör konstprojekt.
En äldre man springer på en livlig gata.
En rödhårig flicka som ler bredvid en brunhårig man som också ler.
Barn ber innan skolan börjar.
En kvinna i vitt och en kvinna i svart står bredvid varandra och pratar på mobiler.
En kvinna och ett barn sitter tillsammans och ler.
En kvinna med svart kjol och pumpar rider sin vita och röda moped.
En grupp av flera personer som står runt ett räcke
Ett rött tvåplan på himlen, med ett spår av rök.
En afrikansk kvinna skakar damm ur något.
En hockeyspelare ligger på isen framför målet.
En person på en bmx cykel, kör en kurs.
En stor grupp människor går nerför en gata, en del bär flaggor eller banderoller.
En kvinna använder en symaskin som barnklocka.
Två skateboardåkare, en med svart t-shirt och den andra med vit t-shirt, tävlar mot varandra.
Flera människor pratar i en gränd.
Childern leker på en karusell som vuxna på en bänk tittar på dem.
Två bergsbestigare nära basen av ett rockansikte.
Många människor sitter vid långa bord fyllda med datorer men de flesta använder dem inte.
En ung kvinna hoppar på en studsmatta
En pojke på en skateboard balanserar på en röd stråle.
En man i blå uniform sparkar fotbollen nerför planen
En person i en vit skjorta som skateboardar på en räls.
Två hundar springer tillsammans genom klippt gräs.
Skateboardåkaren är på väg att hoppa från en träbänk.
Två barn spelar fotboll tillsammans.
En man i brun hatt står upp i en grupp.
Äldre man som sätter på strumpor i en trädlös sanddyn.
En arbetare förbereder fisk för försäljning på en marknad.
Blond flicka i grön klänning med rosa blommor.
Tre ballerinor klädda i vitt, dansar utomhus medan en kvinna i svart klänning ser på.
En blå buss står parkerad på gatan, en man går förbi.
En man i grön hatt och blå badbyxor solar på stranden.
En man som läser en tidning på soffan.
Det finns tre kvinnor i olika klänningar och pannband som dansar på gatan.
En cyklist förbereder sig för att gå nerför en kulle.
En gråhårig kvinna i en grå halsduk och en svart skjorta sitter ett bord med en plastpåse i handen.
En person sover på trottoaren med sitt ansikte täckt.
En kvinna med namnet Steph på sin gula skjorta deltar i ett löplopp med andra racerförare.
En kvinna med solglasögon går på trottoaren.
Många människor samlas runt en gata med träd som talar.
Gondolen rullar sin båt i kanalen.
En man som knäböjer på marken omgiven av flera katter
En kvinna poserar bredvid ett snurrande hjul.
En man är på väg att tacklas i rugby spelet.
Flera människor kör ett lopp bredvid en vingård.
En baseballspelare håller sitt slagträ, medan catcher och umpire huk bakom honom och en publik tittar.
En liten pojke springer över en korsning.
En ensam segelbåt rör sig över ett vackert blått hav med två man vid rodret.
Två män med fiskeredskap pratar utanför.
En kille flyger genom luften på sin cykel i en skateboardpark.
En kvinna sitter på ett tåg och läser uppmärksamt.
En skateboardåkare högt uppe i luften ovanför en inomhusramp.
Den bruna hunden springer ut på gräset.
En vit hund jagar ett uppstoppat djur som dras i ett snöre.
En hund hoppar på trottoaren.
En löpare med rutiga shorts kör ett lopp på landsbygden.
En grupp människor springer uppför en kulle.
Runners deltar i ett lopp kör upp en kulle på en asfalterad väg genom vinlandet.
Två män utför dagliga uppgifter på en livsmedelsmarknad.
En person tumlar på marken bredvid en annan person med skorna av.
En kvinna som dyker i en blå baddräkt.
En man med vita skor, en vit hatt och en vit skjorta som springer på trottoaren.
Män och kvinnor bär rött på gatan.
En snowboardåkare i luften över ett snöigt berg.
Två hundar leker på ett gräsfält
En kvinna står på en bro med en folkmassa bakom sig.
En man som rider på en häst och hoppar över ett trästaket.
Folk som sitter vid ett picknickbord i ett gräsområde nära ett träd.
Fyra personer dansar på en öppen gata.
Två hundar på gräset som skäller på varandra.
En brun hund och en svart hund som leker med en gul fotboll.
En man som spelade cricket pekade mot himlen.
En häst och ryttare hoppar ett litet staket.
En man i långärmad skjorta som rider en gul moped tvärs över en gata.
En pianist och en sångare är redo att uppträda.
En kvinna i svart sitter bredvid en man som bär glasögon i ett kafé.
En man i blått fångas direkt efter att ha släppt bowlingbollen.
Två husky små pojkar i svart klänning skjortor med långklippta frisyrer står bakom den sittande kvinnan i den vita blusen.
En man som gör krattan till sin bästa vän.
En man hoppar på en grön cykel över en skylt som säger "fri middag".
En person som fotograferar ett barn i färgstarka kläder.
En brud och brudgum står tillsammans framför ett trästaket.
En hund fångar en boll i luften
En brun hund hoppar i luften för att fånga en vit volleyboll.
Två män slåss i en boxningsmatch med vita handskar.
Två män boxas i en match.
En man som kikar ut genom ett fönster i ett handelshus.
En grupp barn leker runt i vatten.
Två boxare med vita handskar slåss.
En hund med en repleksak i munnen springer på gräset.
Män som uppträder inför en folkmassa.
Flera barn står runt på gatorna en leker med en boll
Ett par gifter sig, bruden håller rosa blommor.
En person simmar i en vattenförekomst med ett vattenfall.
En gammal flintskallig man i rampljuset som spelar gitarr.
En sittande man som spelar en liten gitarr bredvid en stående man som plockar en bas.
En man i cykelhjälm pratar på en mobiltelefon med andra bakom sig.
Tre män sätter sig ner i en byggnad upplyst med grönt ljus.
Två flickor och en pojke dansar.
Vuxna och barn leker med vattenballonger på gatan.
En grupp människor som står på gatan
En löpare gör ett ansikte under ett lopp eftersom han har ont.
Folk sitter på byggnadsställningar på en stor, vit byggnad.
En ung pojke i röd uniform hoppar på en studsmatta.
En kvinna och en man i tröja instruerar många små barn inomhus
En grupp asiatiska barn spelar ett spel genom att stå i en cirkel bland andra vuxna.
Asiatisk ung pojke med en grå tröja, spelar en asiatisk spel.
En person som bär en grå och röd jacka som löper genom sanden mot bergen.
Flera vuxna pratar med en grupp barn.
En grupp människor går nerför en stig i ett skogsområde.
En far och son tar en paus.
En kvinna och ett barn, både med mörkt hår och ögon leker med två valpar som ligger på marken.
En man som ler medan han håller en akustisk gitarr.
En man som bär en gul hjälm klättrar upp på sidan av en stor stenvägg.
En liten båt som bär två personer rör sig genom vattnet.
En man plockar upp och svingar ett litet barn medan ett annat barn ser på.
En liten flicka som blåser en bubbla bland andra barn.
Två asiatiska män leder en grupp barn i ett spel som innebär att röra ditt huvud.
Två barn läste i sängen.
En svart och vit hund simmar i lite vatten
Flickan är i parken och leker på djungelgym.
En ung pojke som bär hjälm och cyklar i en park.
Man kysser en kvinnas nacke på en livlig trottoar.
Två män pratar vid en tegelvägg.
En person bakom några väskor inuti en igloo.
En man åker nerför en snöig kulle med ett stort berg i bakgrunden.
En man sitter och spelar sitt instrument när parkbesökare sitter bakom honom.
Fyra personer sitter på en stenmur med utsikt över träd och byggnader.
En flicka hoppar ett hinder och kommer att röra marken.
En gammal kvinna sitter bredvid en ung flicka med fingrarna i munnen.
En barfota man på en kulle är böjd över.
En man som ska kasta en leksak för en hund att gå och hämta.
En byggnadsarbetare, mitt på gatan.
Lång svart man står med en hund i förgrunden, en annan svart man i bakgrunden tittar över scenen.
En man sitter på en bänk och lagar mat.
Två män arbetar på kloakerna mitt i vägen som en BMW stannar bredvid dem.
En blond kvinna i en brun skjorta som skickade ett sms.
En inline åkare i röda byxor och blå skjorta skridskor mellan gröna kottar.
Sportspelare öppnar en flaska champagne för att fira sin seger
Mammahunden matar sina ungar.
En närbild av en kolibri.
En motocross ryttare reser längs en grusväg med människor som tittar.
3 tjejer har kul när de spelar kortspel.
En kvinna går med sin son som har en ryggsäck med koppel.
En hytt skott av ett mycket trångt flygplan
En flicka är i luften med kablar bundna till henne omgiven av blå himmel.
Ett par har en diskussion på kanten av en kanal.
En basebollspelare, i vit uniform och röd hatt, gör sig redo att kasta en boll på en solig dag.
Två män som uppträder rör sig nära havet.
Den stora vita fågeln sveper ner svävande ovanför vattnet.
Den svarta hunden rinner genom vatten.
En man sitter ute på ett trästaket mitt i ett stort gräsfält i morgonsolen.
Två personer en man och kvinna rider en elefant på ett fält.
Tre elefanter, som var och en bär på en grupp människor, går genom vattnet.
En man spelar gitarr på en trottoar medan det regnar.
En man dricker på en drink medan han lyssnar på en gentleman som pratar med honom.
Två män springer genom en parkeringsplats med kamouflagebyxor.
En kille som mal över en kant i sin skateboard.
En gymnast gör ett handstöd på de parallella barerna.
En studentmusikensemble repar ett stycke musik.
En ung flicka kastar upp sin examensmössa i luften.
Två svarta hundar leker med en orange stoppad hundleksak.
En flicka står på en snöig klippa.
Ung pojke med brunt hår och svart goggles koppande händer över ansiktet som växer fram ur vattnet i en pool
Flera personer på en buss, en är en olycklig kvinna.
Man med gevär, glasögon, hatt, i kamouflage tar bilder bredvid hund, framför ett fält.
En musiker och en publik bredvid scenen full av musikinstrument.
Två unga pojkar leker i vattnet.
Tjej i rosa toppdans på ett fält.
Kvinna med röd hjälm och röda och svarta strumpor spelar roller derby.
En man som åker vattenskidor genom luften nära en docka.
En flicka i cowboyhatt och en pojke som står på havets strand
En man jobbar i en cykelaffär.
Ett barn i en vit och grön fotbollsuniform sparkar en vit boll.
En liten pojke med orange skjorta sitter på en lila stol.
En kvinna som åker skridskor i en roller derby med en röd hjälm med en vit stjärna på.
Ett asiatiskt barn är naken och har kul i vattnet, trots att det ligger i smutsigt vatten.
En vit och solbränd hund löper längs det gröna gräset.
Två män spelar lacrosse eller fälthockey.
Tre pojkar i kostym, sashes och en flicka i en klänning i sash på ett fält.
En fyrhjuling skickar jord som flyger upp i luften.
Tre män i svarta jackor står vid ett skrivbord i ett fält som håller röda mikrofoner.
En grupp barn sitter, står och knäböjer längs en vägg.
En man i ett resecentrum bär på många saker.
Det lilla barnet står på en trehjuling.
En man i en röd uniform svänger medan en annan i en blå uniform hoppar och andra tittar på.
En skateboardåkare närmar sig en ramp.
Personen kastar ett gult föremål i luften medan han står på sanden.
Ett barn med röd kort på väg att hoppa in i poolen
En grupp löpare som står framför en röd bil i Europa.
De två männen är engagerade i en boxningsmatch.
Tre personer går genom ett skogsområde under dagen.
En kvinna som städar en nysskärm på en restaurang.
En brun hund står på bakbenen och försöker nå något i mannens hand.
En person som hoppar en ramp med tre personer i bakgrunden.
Två kvinnor i svart med flaggor står framför en gammaldags bil.
De tre männen spelar basket på en blacktop.
Tre personer hukar sig ner nära marken med orange hinkar bredvid sig.
En kvinna lämnar tillbaka tennisbollen.
En man i brun rock och jeans går nerför en gata.
En man i en grupp människor tar ett foto.
En röd racerbil som kör på en grusväg med en grupp människor som tittar.
Det blå och grå fordonet är racing genom gruset.
Cyklist rida kursen nära havet som dagen kommer till ett slut.
En man på en cykel gör ett mycket högt hopp.
Det här är ett gäng människor som står i kö vid vad som ser ut som en cykelaffär.
Man i brun skjorta matlagning kött matlagning kött på en liten grill.
En brun hund med en blå munkorg springer på grönt gräs.
Tre unga män inspekterar sina cyklar i solen.
En rad cyklar, och människor som sitter på en brygga, nära vattensidan.
Vissa är i en cykelaffär.
En kvinna i en grön topp som cyklar.
Individuell på klippor med ett vattenfall i bakgrunden.
En ung pojke som bär kostym och hatt håller hand med en flicka i grön klänning.
En person som skateboardar nerför en ramp på natten.
Fyra musiker står och spelar sitt instrument och sjunger in i mikrofoner.
Två personer i flytvästar i en roddbåt
En stor grupp människor tittar på något, skriker och tar bilder.
En sjabbig man står nära en vagn full av lådor.
En ung pojke med röd skjorta, blå jeans och sneakers tycks löpa förbi Pioneer Countys kontor.
Flera människor klättrar upp i ett snötäckt berg.
Två vita svanar i sjön.
En nybörjare gymnast visar hennes akrobatiska talang genom att hoppa från en bar pall.
Män i uniform, med flaggor, samlas utomhus för en ceremoni.
Nummer 24 tycker att det är hans tur att göra mål fotboll.
7 personer som bär alla svarta går på en glaciär.
En kastare kastar bollen.
En kvinna klädd i blått hoppar in i vattenbrynet vid en strand när en fotograf tar en bild.
Turister står en bergsvy under en klarblå himmel.
Två personer med röda västar står i vit snö i en passage.
En nascar förare försöker hålla sin bil på banan
En hund som springer på stranden med en man som tittar i bakgrunden.
En pojke står på en svart bänk.
En pojke i grönt kastar sitt vänstra ben i en spark.
Tre svarta hundar springer efter en orange boll.
En man med hatt och en kvinna med svart topp går på en gräsplan.
En man i gul skjorta håller tummen ute.
Två unga män på cyklar en gör en vända medan den andra klockor
En man i solglasögon som sitter bredvid ett bord fullt av drycker.
En man i den blå skjortan spelar en låt på sin gitarr medan en kvinna och ett barn lyssnar.
Muskulära man tar bilder av en sjö med båtar.
En person cyklar på en grusväg.
Man paddlar röd kajak, orange kajak i bakgrunden.
Två valpar sliter på en trasa i gräset.
En polis på en häst omgiven av åskådare.
En man kastar en frisbee till sin hund som hoppar för att fånga den.
Ett leende litet barn i en rosa baddräkt ligger i vattnet.
En grupp barn hålls samman på en gård med ett bambustaket.
En person i en lång kappa och en käpp som går.
Tre unga män står mot en vägg och pratar medan en ung pojke ser fram emot att hålla en affisch.
En man gör Ti Chi på en klippa med utsikt över en skog.
Två kvinnor och en man är klädda vid ett bord runt en lykta i skogen.
Pojken i den röda skjortan skateboardar.
Två tonårspojkar hoppar in i en hotellpool.
En del människor väntar på att köpa varor från en gatuförsäljare.
Två klättrare bär ryggsäckar som stiger upp i ett mycket snöigt berg.
Två människor klättrar upp för ett stort, snöigt berg.
En tjej i rosa hoppar upp i luften i en bowlinghall.
Två vuxna njuter av en målning av handavtryck.
Tonåringar poserar för en bild på en fullsatt händelse.
En ung flicka i en ljusgul klänning omgiven av gula blommor
Säljaren håller en hel del ballonger som skapats i form av Disney tecken.
En man klättrar upp ur havet på en klippa
En man med akvabyxor och matchande flip-flops drar en vagn med handgjorda kvastar genom gatan.
En man i gul skjorta står vid en disk.
Två kvinnor i en blandning av islamisk och amerikansk dräkt tar med sig stora lådor på en vagn genom en utcheckningslinje.
En asiatisk man som cyklade nerför gatan.
En rad militära lastbilar passerar förbi en soldat som går sin väg.
En kvinna som sätter ett halsband på en annan kvinna
En fågel flyger ner till marken.
En hund som plaskar genom en pöl i gräset.
Två kvinnor som bär hjälm och skyddskuddar verkar slåss.
En kvinna i rosa jacka sitter medan hon skriver på en laptop.
Pojken i de svarta badbyxorna dyker ner i poolen.
En dykare under vattnet poserar bredvid en stor akvatisk organism.
En liten pojke i vit skjorta hoppar med ett svärd i handen.
Man i kampsport stil kostym hoppa i luften.
En fullsatt buss och en ung man i glasögon som nyper näsan.
En person som lär sig att klättra med en annan person hjälper till.
Två män klättrar på en intressant formad klippa.
Tre personer, två spela trummor och en spela ett horn instrument.
En cowboy vinkar en lasso i luften på en hästshow.
Tre poliser, en på poliscykeln, bär svarta uniformer med svarta stövlar.
Gatuutsikt över en stad med en gammal asiatisk kvinna som går förbi en telefonkiosk.
Två unga barn går uppför några trappor.
En brun hund trampar vattnet med något i munnen.
Två personer stannar på en tom stad gata.
En person cyklar med en röd vägg i bakgrunden.
En fläckig svart och vit hund stänker i vattnet.
Två flickor poserar bakom ett träd med stora leenden.
En grupp barn åker tunnelbana.
En pojke som gör en volt i luften på stranden.
En svart hund sticker näsan i vattnet.
Fyra unga kvinnor i bikini baddräkt hoppar ut i havet en solig dag.
Peoople står utanför en byggnad nära en gata.
Folk på gatan tittar på en gatuartist med gitarr.
En brun hund hoppar i havet.
En grupp människor rider hästar genom ett skogsområde.
Damer som tas genom en övning rutin av militären
En man klättrar upp på en klippavsats.
En pojke klättrar upp i ett träd och ler för bilden.
Tre flickor i färgglada kläder dansar under ett scenljus.
Två män och en kvinna som spelar ett lyckligt spel av snurra flaskan.
En amerikansk armésoldat lär en student hur man behandlar sår
En grupp vuxna har sina cyklar redo att rida
En soldat som går en hund med en väska i munnen.
En kvinna skriver på pappersarbete vid ett evenemang.
En flicka gör en sidoböj i surfingen, en annan flicka bakom henne, solen går ner.
Tre personer lastar eller lastar av sin bil.
En kvinna bär ett barn över en stenbro.
En mycket glad person som går i skogen med löven blåser.
En ung flicka upp och ner på en swing set
En kvinna står framför en man som håller ett litet leende barn.
En baseman fångar en baseball medan en löpare glider för att röra vid basen under ett basebollspel.
En fastare rakning utanför medan en hund är vid hans sida.
De flesta sitter vid bord och läser, men en man ser ut att sova.
En man och kvinnor arbetar med varandra
En liten skara människor som sitter vid bord och äter mat eller dryck medan andra står eller går.
Den Red Sox outfielder fångar en fluga baseball med sin handske.
New York Mets avslutade inningen genom att fånga en alltför ivrig Boston spelare på väg tillbaka till första.
En grupp människor lyssnar på någon som pratar.
Två hundar springer med ett litet barn längs en sjö
Kvinnor som sitter i stolar tittar genom ett bindemedel.
En man kör motorcykel i smutsen nära buskarna.
En man i blått som hoppar på en smutscykel.
En kvinna som bär en uppvärmningsdräkt tittar på sin mobiltelefon.
En ung hona med brunt hår håller en orange fjäril.
En grupp män sitter och står på en gård, en del läser böcker och en del pratar.
En flicka klädd i rosa springer från havet till stranden.
Två unga män och en kvinna står på baksidan av en blå pickup som sorterar genom grönsaker med leenden i ansiktet.
Tjejen i rosa randiga vantar skrattar i folkmassan.
När man sitter på en blå plaststol, skalar en man i rosa skjorta frukten i en skål.
Ett köp skateboard på en skateboardpark.
Mannen utför ett trick på en motorcykel högt i luften.
En brottare hoppar över repen.
Två personer tittar ut i vattnet i slutet av en träbrygga.
En blå fågel flyger genom träden.
En man som dricker ur två gröna vinflaskor samtidigt.
Ett barn i svart skjorta tuggar en blå elefantleksak.
Spädbarnspojke med blont hår i blå täppa sandaler, blå hoppare, vidrörande en orange trafikkon.
Ett barn som ritar en bild med kritor
Två racerbilar på en väg framför en gräsbevuxen parkeringsplats.
En man och en kvinna som tränar i en park.
En stor kvinna i en svart och vit rand skjorta håller några färgglada dekorationer medan stirrar på två män.
En liten pojke i en grön randig skjorta som håller upp en pinne på verandan.
En grupp människor som ler och rider på en båt.
Mannen bär flera lådor medan han åker skateboard.
En man åker rullskridskor nerför väggen bredvid några vita trappsteg.
Par sover på tunnelbanan bredvid varandra.
En man sover på en bänk bakom en fontän.
En ung pojke i patriotiska shorts som springer på stranden.
En leende blond-hövdad liten flicka ligger på golvet magen ner tittar upp medan en rad dominos sitter bredvid henne.
En pojke och en flicka kysser varandra i solnedgången.
Två hundar, en solbränna och en svart, leker dragkamp på gräset nära dammen.
Barnet tycker om att bada.
Två asiatiska kvinnor med kort svart hår som pratar med varandra.
Många människor sitter ett bord klädda bord äta mat och göra samtal.
Hane i grön rutig skjorta och namnskylt, håller en mikrofon med höger tumme i sin blå jeans ficka.
En man i grön jacka som röker en cigarett kastar en liten boll.
En kvinna pratar med sina vänner när hon sitter på en restaurang.
En ung pojke simmar med glasögon.
Flera kvinnor klädda i zigenarliknande kläder dansar omkring i en skog.
En hund går på en stig omgiven av träd.
En kvinna som bär en gul skjorta löper längs ett rött spår.
En man interagerar med en hund som springer förbi honom.
Det finns män i ett rum med läsk och chips på ett bord.
Man spelar ett spel med en ung flicka.
En liten pojke med glasögon håller i en pistol.
Tre kvinnor i affärskläder går över en gårdsplan.
En kvinna sitter på en buss mot många bruna hus.
En flicka ligger på en kort tegelvägg.
En brindlehund som står bredvid ett julgransträd och sniffar ett litet barn som ligger på golvet när barnet leker med leksaksfordon.
Ett barn i rosa klänning utanför.
En ung flicka i gul klänning och en liten pojke i vit kostym.
Vattenskidåkare hoppar från vattnets yta, okänd struktur i bakgrunden.
En man som står bredvid en liten flicka som står i en soptunna på en gård.
En gul hund springer genom grönt gräs.
Två tonårskillar gör skateboardtrick på en skatepark.
Mannen och barnet simmar.
En man hoppar från en klippa ner i havet medan andra tittar.
En man i nyanser och en tröja ser en flicka stå i en återvinningsbehållare.
Pojken som bär den röda jackan hänger på sidan av gungan.
En ung dam bär ljusrosa solglasögon och sitter på en liten studsmatta.
5 manliga polospelare i aktion under ett spel på en poloplan på en solig dag.
Två kvinnor klättrar över klippor nära havet.
Två pojkar går ut på ett militärmonument över gräsiga gröna fält.
De tre hundarna leker i sanden.
Sex personer poserar för en bild framför en vägg med graffiti.
En kvinna som bär hjälm är i en rullskridskotävling.
En man med rakat huvud står i en flod och håller i ett rep.
Två brindle hundar springer i gräset.
En kvinna i svart och blå kläder dansar på gatan med en kvinna i svart och röd utstyrsel.
En man som grillar korv och korv.
En baseboll kanna i en röd och vit uniform kastar bollen medan hans lagkamrat tittar.
En kvinna i en orange halsduk drar ett paket cigaretter ur en kartong.
En publikscen med människor i gula och vita infödda kläder.
Vuxna som bär ballonghattar ser barn leka i ett ballongslott.
En jockey rider på en kurs.
Äldre par dansar på natten, med ljussträngar i bakgrunden.
En ung pojke i en grön gunga rider genom luften nära en lada.
En man sitter vid sjön, under ett paraply och målar.
En flock måsar lyfter från stranden.
Två pojkar gunga stående upp på en gul gunga uppsättning
Tre mountain bikeers är i ett lopp i skogen.
En grupp pojkar spelar basket tillsammans.
Ett blått, rött och gult plan gör en slinga i luften.
En ung pojke som tar en bild genom glaset och två honor som pratar.
En vit hund och en svart och vit hund leker medan ytterligare två svarta hundar rör sig mot dem.
En man som sitter i en stol framför en röd byggnad.
Två kvinnor, som är mycket atletiska, spelar beachvolleyboll.
Person som gör en skateboard stunt
Fyra unga valpar kramas ihop mitt i en filt.
Tre valpar ligger på en soffa bredvid en barnflaska.
Två vita och bruna hundar skäller på strandlinjen medan vågorna rullar in bakom dem.
Två vita hundar och en ljusbrun hund som springer längs stranden.
Två kvinnor visar olika ansiktsuttryck och bär guld och lila kostymer.
En flicka som leker i en pöl när hon bär en rosa rock
Fadern och en son springer i havsstranden.
En man med svart hatt som öppnar en kartong.
Två pojkar sparkar en gul fotboll i surfingen på stranden.
En man med ljusblå skjorta och marinbyxor går nerför en gränd.
En hund simmar genom djupt vatten nära flera ankor.
Två män sparkar.
En man tittar över en meny medan servitören väntar på sin beställning.
En varmluftsballong har svårt att lyfta.
Flera små barn med fingertopparna på en vit frisbee
En äldre man i en vit tröja pratar på en mobiltelefon.
En man klädd i en orangefärgad rock klädd i sandaler sitter på en bänk utanför en byggnad.
En grupp barn och en mamma tittar på när en amerikansk flicka spelar på sin mobiltelefon.
Två barn skrattar och leker i en däcksvinge i en park.
Ett litet barn som sitter på knä på ett vitt kakelgolv.
En smet svänger på en baseball med en smet som värms upp i bakgrunden.
En liten pojke som slåss i en basebollmatch.
En person som tar en bild av någon som åker skridskor ner för ett räcke på natten.
En anka flaxar sina vingar nära vattnet.
Tre byggarbetare som tar en paus i närheten av sin fabrik.
Den brunhåriga mannen och kvinnan poserar för en bild.
Det finns en person som står i vatten och leker med en hund.
En indianhövding i full klänning.
Ett amerikanskt band spelar instrument under ett tält.
En ung man med en brun skjorta som hoppar högt i luften på mattor.
Folk tittar på två män i brungula dräkter som hanterar ormar på grusväg.
En ung man hoppar en cykel från en sluttande vägg över en bänk.
En man utan tröja gör ett trick på sin röda och svarta cykel.
Två motorcykelförare på ett spår, en utan sin motorcykel.
En grupp kvinnor som rider på hästar medan de håller flaggor från flera nationer
Tre personer brottas med en tjur på en rodeo.
En kvinna med gitarr sjunger framför en byggnad och gräs.
Tre personer står på promenad och tittar på byggnader tvärs över vattnet.
En labbhund står på en fallen trädstam med en kille i bakgrunden.
En kvinna i en blå tennis outfit avslutar en swing.
En man med lila hatt och clownmakeup hejar på folk.
En man på en rodeo kastas av en häst.
En kvinna får sitt hår hoprullat av någon annan med locktång.
Män på rodeo försöker tämja en tjur.
Mannen i svart flyger iväg framför ett rött staket.
En hund hoppar genom ett snöigt fält.
En kvinna hoppar upp för att undvika en läcka från en jäsningstank.
Ung pojke med röda badbyxor som leker i sand på stranden.
En kille med blå hjälm står på rep ovanför alla andra.
Man spelar gitarr i ett mörkt rum.
En man med en käpp i vänster hand på ett fält
En cykelcyklist rider i motsatt riktning av trafiken.
En man går över ett tak i staden med en drake som flyger ovanför.
En man som ramlade av sin surfbräda.
En surfare på en gul surfbräda stänker upp vatten på en annan surfare.
Man sätter upp bord med osthjul.
En grupp hockeyspelare och en officiell monter på isen under ett spel.
En kvinna som går parallellt med en gul linje mot trafiken.
En kvinna arbetar i en monter med färgglada varor.
Örnen flyger ner till marken.
Två kvinnor dricker och roar sig.
Man paddlar förlora sin paddel och faller ur båten.
En man med rakat huvud på mountainbike.
En liten svart hund hoppar över en bar.
En man och en kvinna som håller muggar med en annan man i närheten.
En stor grupp människor vid sammankomsten av något slag som använder sig av varor.
Gul hund står på bakben med boll i munnen, bygga i bakgrunden.
Två kvinnor sitter vid ett bord och arbetar tillsammans med hantverk.
En ung flicka som gör ett konsthantverksprojekt som lärare tittar över bordet.
En äldre kvinna skär något ur en bok.
En del lärare gör pyssel och de andra diskuterar något i ett färgglatt rum.
En grupp kvinnor som dansar tillsammans.
En brun hund springer på en sten.
Barn spelar fotboll, medan en vuxen tittar på.
En ung kvinna med tajta magmuskler lyfter vikter.
Två personer äter mat i solljuset.
En man utan skjorta och ryggsäck har en låda på huvudet.
Åskådare som tittar på en motorcyklist marken runt ett spår.
Det finns ett träd eller en vinstock på sidan av byggnaden.
Männen använder horor för att bryta jorden.
En pojke gör ett skateboard trick i luften.
En pojke med en basketboll som hoppar mot målet.
En flickas händer, en annans fötter och en pojke som spelar bongofat sitter på ett picknickbord.
De två pojkarna leker i våt sand.
Den unga kvinnan med scarfen ger en present till någon.
Killar samlades utanför en glassaffär en solig dag.
En brun och vit hund springer i ett fält av gula blommor.
En grupp människor har fest.
En grupp personer med bagagelinje utanför en flygplats.
En svart hund som går längs en stenig terräng.
Dottern medger att hennes mamma är cool i sina flygarsolglasögon.
Två asiatiska kvinnor har en livlig YMCA-affisch.
En man i grön kajak paddlar genom vattnet.
En pojke som slår med en snösprej.
En kille får håret avrakat av en annan kille, medan en tredje tar en bild.
Fyra barn väntar som någon skär trä.
En man som bär ryggsäck tittar upp mot ett vattenfall.
En hund som springer på en stig i bergen.
En man i grå skjorta viftar mitt i en plantskola
Mamma och barn med blå skjortor som leker utomhus.
En skateboardåkare gör ett trick när det gäller att hantera en skål.
Folk går på en trottoar i en stad.
Tjejen gör en konstig ansiktsdans i en parad.
En jockey som svider en häst förbereder sig för att hoppa över ett hinder
En kvinna som bär en svartvit dräkt är skickligt isåkning medan andra tittar på henne.
Två barn i blå skjortor som ligger på bänkar
En kvinna i solglasögon ler när hon sitter ovanpå några stenar.
Två män i olika färgade tröjor spelar hockey.
En man är delvis silhuetterad och lutar sig mot ett mörkt föremål.
Jockeys på hästar under ett lopp.
En man och en kvinna som kysser inför en massa människor.
Röd och vit motorcykel nummer 58 tävlingar runt banan.
Två män står nära en metallkonstruktion framför en tegelvägg.
En unge som rör en baseball och bär en blå hjälm.
En pojke med en t-shirt på som säger FROG! står blad genom sidorna i en bok.
En man på en cykel utför ett hopp.
Två män i skyddsvästar arbetar med ett projekt utomhus.
En gata med flera personer och flera handelsbodar längs båda sidor.
En liten svart hund i havet med några stenar i bakgrunden
Två byggnadsarbetare slätar ut betongytan.
En liten flicka står bredvid en annan liten flicka som tar ett fotografi.
Baseballspelaren är ute efter bollen.
En man i orange hård hatt som använder tunga maskiner.
En grupp män som spelar Lacrosse på natten.
Dansare i vitt uppträder på en mörklagd scen med en rosa upplyst nyans som lyser upp dem.
En våt hund som leker med en leksak i vattnet.
En pojke kastar ett föremål i luften medan några andra barn tittar på honom.
Racing på våt väg medan människan hänger på baksidan.
Mannen ser väldigt spännande ut med hörlurarna stående utanför bredvid en kvinna.
En grupp människor som dansar tillsammans.
En kvinna i blått och en man i rött är på väg att kyssas med lövverk i närheten.
En man, som låg på gräset, räckte ut handen mot en annan arm.
En man klädd i blått stående framför en färgglad frukt- och grönsaksställning
Cheerleaders, bygga en pyramid, posera framför en publik.
Två hejaklacksledare klädda i svart och rosa poserar med ett ben som hålls upp.
Cheerleaders i Falcons kläder bildar en pyramid.
Två personer och en hund leker i vattnet med hjälp av en blå uppblåsbar leksak.
Ung flicka i röd klänning kysser en annan tjej på huvudet.
En grupp barn samlas runt en vit hund på gräset utanför.
Ungdomar sitter och pratar i en kaffebar.
Den stora hunden tittar genom staketet på den lilla hunden.
Mannen inspekterar sin cykel nära en väg.
En liten pojke med blå skjorta bär en blå spade på stranden, när han springer mot ett par måsar.
En baseballspelare passerar bollen, medan en man går över kamerans sikt.
Två barn ligger i en pool med en strandboll flytande i närheten.
En grupp hejaklacksledare hejar på.
Det finns en grupp på åtta personer som paddlar kajaker i en vattenförekomst.
En mountainbike racer hoppar sin cykel som åskådare klocka.
Två män i en orange båt rider över vattnet.
En pojke och en flicka leker på golvet med ett tågsätt.
En man i röda badbyxor som knuffar en barnvagn nerför en fullsatt strand.
Två män går framför en vit tegelbyggnad.
En man med blå skjorta spelar trummor.
En man på en skateboard medan publiken tittar.
En silverbil går utom kontroll på en kapplöpningsbana.
En simmare som gör bröstsim i en pool.
En hund står på bakbenen med sina tassar utsträckta medan han bär ett rött föremål i munnen.
Tre nosade och numrerade hundar som sprang genom gräset.
En grupp människor, många med ryggsäckar, går nerför en korridor med rullande bagage.
En man i svart skjorta och bruna shorts äter.
En ung man skateboard i svarta skor, svarta byxor och en vit topp med solglasögon.
En kvinna som spelar på en överdimensionerad checkerbräda.
En tatuerad man med en vit hund som hoppar upp för en pinne.
Två personer på en bänk sitter i skuggan.
Två män som bär hjälm är knäböjda bland sex trafikkottar på gatan.
En man klättrar på klippor vid vattnet.
Två hundar leker i en flod, en gör ett stänk.
Tre barn leker med bollar på en gräsmatta
Två personer utför en dans med eld som huvudattraktion.
En man har två valpar.
En smutscykelcyklist tar en okonventionell stig i ett stenigt område.
En grupp människor rider i en buss.
Ett barn som är under 10 år är mitt uppe i luften under en basketboll.
En ung man sover på jobbet på en stol utanför dörren.
Två barn, en klädd i vitt, klädd i rött, lekte i vattnet på en strand.
Ett barn kastas i luften på stranden.
Nummer åtta rullskridskor tar ledningen och drar sig undan från sina svarta och röda klädda motståndare.
En man ligger i ett litet flerfärgstält.
En grupp människor sitter på trappan utanför.
En man på avstånd som fyller en hjulpipa.
En ung pojke som bär en stor fotbollsboll med en fotboll i bakgrunden
Pojken spelar baseball på ett gräsfält.
En brunett finns utanför en frukt- och grönsaksbutik och väljer matvaror att köpa.
Den stora hunden ser den lilla leka med rep.
Tre män justerar rep runt ett brunt metallrör.
En hund vadar i vattnet
En man hoppar med kroppen framåt mot en fotoskärm och ett stort fotoljus.
Barn i uniform går till skolan.
En man i grått sitter och tittar på ett vattenfall från en klippa.
En grupp som arbetar tillsammans för att dra något åt land.
En vandrare passerar en vit klippformation mitt i en tom öken.
En ung pojke i en blå transformatorskjorta som går i grunt vatten med en glad look i ansiktet.
Ryttare på en berg- och dalbana håller händerna uppe i spänning när tåget springer nerför spåren.
Den unge mannen hoppar för att servera volleybollen på stranden.
Två män i en bur boxas med varandra inför massor av människor.
Tre personer rider på en blå och vit båt.
En pojke i vit skjorta gör en spark i luften.
En ung man i en fiskekanot.
En ung pojke som bär en spindelmönsterskjorta på sanden.
Damerna med den här unga flickan ser lyckliga ut.
En man är på baksidan av sin vän.
Två män hoppar runt tillsammans utanför en byggnad.
En pojke ryggar tillbaka från sanden på sitt blotta bröst.
En man som maler ner en ledstång.
En blond kvinna i en grön tank topp rider sin cykel framför en lägenhet byggnad.
En professionell brottare hoppar på en annan utanför ringen.
En grupp spelare jagar en boll på ett fält.
Det leende barnet har bubblor nära örat.
Fyra personer går nerför gatan och en försöker hoppa i en kundvagn.
En hund simmar i vattnet.
Pojken på en skateboard hoppar genom luften.
En motocross förare hastigheter av under ett lopp.
En grupp kvinnor i infödda kläder sitter på golvet.
Ett par svarta hundar springer i surfingen.
En man gör ett skridskot trick från graffitifyllda trappor.
Kvinnan i en blå jacka sitter vid kanten av en tennisbana.
En brun och vit hund springer med munnen öppen över ett fält.
Ett fotbollslag poserar för en bild.
En del människor står runt en stor uppblåsbar rutschbana och ser ett barn glida ner för den.
En kvinna med digital klocka sjunger in i en mikrofon.
En mycket glad pojke klättrar upp på en stolpe på en veranda på en bakgård.
Män går med en flock hundar.
Här har vi en kille som använder en trycktvätt på trottoaren.
En flicka i svart hatt som håller i en afrikansk amerikansk bebis.
Ett gäng ungar klättrar upp på ett träd och lägger ner det.
En man med en cigarett i munnen leker pool.
Någon åker skidor från toppen av någon typ av byggnad.
Någon i gul hatt sitter bredvid två fiskestolpar.
Ett barn som bär blå hatt och rock tittar upp på en skylt och pekar.
En ryttare på en gruscykel tävlar genom en skog.
Häst jockeys tävlar på hästar i ett lopp.
En ung flicka i en färgstark utstyrsel kikar genom ett trästängsel.
En kvinna med grön skjorta och en kvinna med orange skjorta poserar med utsträckta armar
Två hästar med ryttare, tävla längs banan.
En man och två kvinnor är inne i ett växthus håller trädgårdsverktyg.
En äldre man står på trottoaren och målar utsikten.
Två män sitter vid ett bord på trottoaren under en francisco gatuskylt
En ung man och kvinna kramar när de bär peruker.
En man i en grön jacka som stirrar på himlen nära en forrest.
En äldre man och en yngre man bär jackor.
Två fotgängare passerar en restaurang titta på hunden som tittar på dem.
En svart och vit hund som hoppar över ett hinder.
En ung flicka sitter framför en maskin som trycker på knappar.
Elever som sitter i en föreläsningssal och lyssnar på en föreläsning.
Ett mans- och kvinnopar dansar med suddiga träd i bakgrunden.
En man och en kvinna som bär röd omfamnande.
En man med byxor och en röd skjorta dansar med en kvinna i en tajt röd klänning.
En man går förbi en röd byggnad och bär specialutrustning.
En vit hund hoppar upp ur vattnet för att fånga en tennisboll.
En hund hoppar över ett hinder.
En coach och domare har en diskussion medan en baseballmatch pågår.
En liten flicka som knäböjer på en säng.
En äldre herre och dam som står på en utomhustrappa och pratar, var och en med mappar i sina händer.
En man sitter utanför bredvid ett träd och buskar.
Två barn sover medan de vuxna dansar bort natten.
Man går bredvid en häst som drar en kärra i skogen.
En ung kille som bär allt grått och en mössa tittar på en boxningssäck medan andra tittar på.
En grupp människor tillbringar tid i en park i kostym.
Sex unga vuxna, en som håller en hund i kopplet, hoppar excstatiskt på stranden.
Skateboardåkarna försöker stunta på natten.
En person är i luften på en cykel nära en vattenförekomst.
Man i shorts och blå skjorta matlagning på kolgrill.
En hoppare rensar ett vitt staket på sin häst.
En man som står i snö med ett berg i bakgrunden
En flicka står med båda händerna uppe och tittar på solnedgången och en segelbåt.
En baby i en pool som stänker vatten i luften.
En man med full huvudmask, khakis, och en blå skjorta sitter på en resväska nära orange och vita byggfat och betalar dragspel för fem personer sitter i gröna och vita gräsmatta stolar.
En man på ett tåg med en blå skjorta på.
En långhårig, skäggig ung skateboardåkare gör ett stunt på en skateboardyta.
Två unga pojkar leker på klipporna.
En brun hund med baseball i munnen.
En kvinna knäböjer inför en symaskin.
Orkester spelar för personer i hårda hattar i ett rum med skadat tak
En man och en kvinna som klär upp sig dansar tillsammans utomhus.
Vit hund med krage löper i inhägnad i gräsyta
Barnet i den blå skjortan springer genom sanden.
En brun hund stirrar i fjärran medan den står på torrt gräs.
En kvinna som tittar genom låssmedens fönster.
En man håller ett stort föremål, böjer sig framför många växter.
En man på ett kontor kollar information på sin laptop.
En svartklädd man surfar på en stor blå våg.
En stor grupp ljusklädda dansare som fotograferar.
Två små flickor läser en bok på biblioteket.
Tre män sitter och skrattar.
En rullskridskor utför ett trick på en ramp.
En man hoppar i luften medan himlen surfar.
Människor är på en utomhus shopping basar promenader och tittar på varor.
Två hundar springer genom ett fält.
En man i flanellskjorta står inne i ett ihåligt träd.
En grupp människor sitter på gula stolar och pratar.
En grupp hundar som står i en flod.
En ung vuxen man står med en basketboll på en plan.
Folk som spelar cricket i parken, tallar där bak.
Två bruna hundar springer genom ett fält.
En ung flicka bär lila skjorta och rosa pannband.
Två terrier hoppar efter en tennisboll i en park
Tre kvinnor och en man sjunger sina hjärtan i mikrofonen.
Två män som bär bagage står mitt i fältet av grönt gräs.
En kvinna försöker rida på en liten våg.
Ett barn leker med en utklädd vuxen på en parad.
Ett litet barn håller en gummikyckling suspenderad i luften
En man med blommor springer från två poliser.
Två kvinnor ler bredvid en mikrofon på en scen.
En blond kvinna står bakom en mikrofon.
Två barn, en pojke och en flicka, som går längs en asfalterad väg och håller ett svart paraply.
Folk går genom ett pittoreskt område.
En man spelar gitarr på trottoaren medan en annan man sitter i bakgrunden nära en cykel.
Den svarta hunden pouncing på något på gården.
Två personer på scenen håller en pose, som andra tecken står på bakgrunden.
Man i gul hatt håller upp trofé
En man på en skateboard som hoppar en orange kon.
Dansare uppträder på scenen.
Den svarta hunden drar i ett grönt rep.
Män med hatt går på gatan.
En äldre gentleman i en rutig skjorta och glasögon ler mot kameran.
Folk på en gårdsmarknad.
Tre stora hundar leker i vattnet på stranden.
En kvinna sträcker sig vid havet vid soluppgången.
Tre leende barn svingar i en däcksvinge på en lekplats.
En överviktig flicka håller en stor svart ökenråtta i sina händer.
En kvinna håller upp sin mobiltelefon till en kartong kattungar medan en annan kvinna tittar på dem.
Två hundar delar en leksak i ett fält av vegetation.
En skara människor som sjunger med fyra gröna strobe lampor skiner i bakgrunden.
En ump i svart tittar på en basebollmatch.
En hejaklacksledare klädd i orange och vit dräkt kastas i luften av fyra andra hejaklacksledare på marken.
Kvinnan visar en stor stjärna av David för unga elever.
En liten flicka i rosa skjorta tar en sväng på en t-boll.
Två personer fotograferas bakifrån sittandes på en buss
Vuxen med glasögon matar en nyfödd kattunge med en liten flaska.
En surfare som går genom en våg.
Dirt cyklister färdas en serie hopp.
En fallskärmshoppare flyger genom luften nära en hög byggnad.
Dessa fyra män, två skjorta utan, skyfflar sand.
Ett sportlag är uppställt utanför.
Flera människor rider cyklar med människor i läktare tittar.
En hund i en "superman" skjorta sover på en filt.
En kvinna i ett stycke baddräkt som stänker i vattnet.
En äldre man sitter och flera personer står.
Två unga pojkar sitter bredvid en färsk frukt monter, på en bondemarknad.
3 båtar i vattnet, person i mellersta båten bär en lila skjorta.
En kvinna i svart tank topp och en man i orange skjorta sitter på ryggen till kameran.
En man som spelar bas på scenen.
En ensam bicyklist med hjälm som hoppar på en graffitierad betongramp.
En bulldozer på en strand utan vatten.
En stor brun hund sitter bredvid en liten vit hund i ett fält av långt gräs.
Den kanadensiska biker sponsras av H&amp;R Block rider av.
En kvinna cyklar i ett cykellopp.
En man håller upp en tävlande i ett cykellopp.
Tre barn bär ansiktsfärg och ler.
Ett barn målar med olika färger med hjälp av borstar.
Mannen utför ett trick högt i luften med en cykel.
En man i röd jacka som klättrar i ansiktet.
Tre kvinnor i saris dans nära en stor flagga.
Två personer som leker med en Frisbee.
Fyra pojkar är ute på en lekplats med en grön och gul boll.
De tre landhockeyspelare jagar alla bollen.
Pojke hoppar från skateboarden när den går nerför trappan.
En liten flicka som målar sidwalken vit.
Fyra män tittar på sin båts motor i floden.
En baseball kastas på ett volleybollnät.
En flicka uppträder medan hon är klädd i en grön och vit randig sari.
Gymnast bär en röd outfit och hoppning.
En man som bär glasögon, en vit skjorta och slips, och slacks står vid en säng som har vita kuddar på sig.
Två unga män poserar för kameran.
Två barn och en man går förbi ett dåligt ihopsatt skjul.
Män spelar baseball.
En kvinna i rött, vitt och blått tävlingskläder som cyklar.
En cyklist gör sig redo att starta sitt inomhuslopp.
En kvinna i pälshatt och svart överrock som sätter på sin vänstra sko.
Ett par står nära vid vattenbrynet.
En man som bär en ljusblå tröja sitter vid ett bord framför en budweiserflaska.
Dessa (7) damer fick en utmärkelse och några fick blommor med en man vid behov.
Tonåringarna vilar på en bänk efter sin löpning.
Cykel racers är racing
En man testar en visning av träningscykelutrustning.
Unga cyklister förbereder sig för ett lopp.
Sex tävlingscyklister väntar på att loppet ska börja vid startlinjen.
En grupp cyklister tävlar i en velodrome.
En pojke gör gymnastik i gräset vid den blå speltunneln, när två pojkar står på uteplatsen till ett hus i ranchstil.
Ungar som spelar boll i parken.
Två hästar tittar över ett staket på ett barn som bär en röd tröja.
En grupp människor samlas på en grusväg nära en bil.
En ung man hoppar över en lång stolpe i en skatepark.
En person torkar ut i vattnet.
En grupp elever som ler framför en kamera.
En brun hund som tittar på en brun hund som simmar i en damm.
En pojke svänger på en gungställning.
Två personer spelar golf på en golfbana.
Flickan i rosa topp rider en skateboard längs en vit vägg.
En hund hoppar genom en röd båge
Det finns grupper av människor i gröna eller lila skjortor samlade utanför hålla tecken och lila ballonger.
En kvinna köper saker från mannen i den röda skjortans gårdsförsäljning.
Två kvinnor, en med kamera, sträcker sig ut och rör vid en spegelkula.
En man i halm hatt och overall är med en vän utomhus.
En leende flicka glider ner för en lila slide fot först.
Ungt par bär formella kläder och dansar långsamt på dansgolvet.
Bruden i den vita klänningen är omgiven av brudgummen och brudtärnorna, alla i svart.
Ett ungt par i bröllopskläder poserar för en bild.
En liten liga fotbollsmatch pågår i ett förortsområde.
En man och en kvinna i bröllopskläder ser ut mot vattnet.
En man spelar gitarr när han sitter på läktare framför en sjö.
Två pojkar sitter och äter glass.
En svart hund som springer i grunt vatten på en strand.
Den utstuderade Jesushelgedomen hålls i en parad.
Män i blått bär något på sina axlar följt av ett band.
En vit kvinna med en Panasonic videokamera i en park.
En surfare som bär en svart och grön våtdräkt som rider på en våg.
Skateboardåkaren rider rampen bredvid den mycket stora målningen.
En skateboardare utför stunt på en graffititäckt skateboardramp.
En flicka knäböjer på en gunga i parken.
En mountainbikeer hoppar sin cykel över en stubbe i skogen.
Fyra brudtärnor poserar dramatiskt med brudgummen.
En ung flicka klädd i röd prick outfit leker med leksak.
En kvinna går fyra hundar.
En tjej med fräknar och metallörhängen njuter av körsbär inomhus.
En man vindsurfar i våtdräkt.
Två kvinnor sitter tillbaka för att backa ut ett kontor område.
En person som spelar cricket i en helt grön outfit
En brunettflygvärdinna i röd uniform knuffar en matvagn på flygplanet.
En hund med gul leksak jagas av en annan hund
En svart hund går på stranden nära klipporna.
En röd lastbil kör över en stenig yta.
En afroamerikansk kvinna går nerför gatan medan hon pratar på en mobiltelefon som håller i en svart handväska.
En man som avslutar lite golvarbete med en pensel.
En asiatisk ung kvinna med vit skjorta och svarta byxor håller i en rosa handväska.
En ung pojke spelar på en gunga.
En stor gul hund och en liten vit hund i gräset.
En man står på en stege uppstött mot en tegelbyggnad.
En kvinna och ett barn tar en tupplur i sanden.
Texas basebollspelare fångar bollen på basen medan motståndaren glider.
En man på en båt gör sig redo att dra i sitt nät för att se vad han fångade.
En grupp på fyra domare betygsätter en tävling.
En man i svart, talar i en mikrofon, medan en kvinna skriver.
Fyra personer sitter vid ett bord framför en publik.
En upptäcktsresande i en isgrotta står ovanför ett stort ark mörkblått is.
Tre cowboys tar en tjur vid hornen och brottas med den.
Två män i svarta kostymer går mot ett kontor.
Någon böjde sig lite i mitten av en stor byggnad.
En man i vit skjorta och en svart keps som sträcker sig upp till en skylt på en tegelvägg.
En man i blå skjorta cyklar på en asfalterad väg.
En blond tjej och brunett brun hängande med gymnastiska rep
En fiskare i en hatt som samlar sina nät i grumligt vatten nära stranden.
En grupp människor som går i samma riktning är två kvinnor, varav en bär solglasögon och shorts.
En ung man som bar en rutig skjorta vid ett tjurslagsmål.
En flicka hoppar från ett högt dyk i en urban miljö.
Asiatiska kvinnor på en fest pratar vid väggen.
Den här skateboardåkaren flyger högt och gör ett trick för att imponera på sin vän.
Ett 5-personsband uppträder på en scen inne i ett tält.
En ung flicka i riddräkt sitter på en häst med en nallebjörn.
En man går ut med två hundar.
Kvinnor i en grön klänning med en lila hulahoop runt henne, en stor skara människor bakom henne.
En man i röd rock är snöblossande på en parkeringsplats.
En liten asiatisk pojke i svart och blå t-shirt står på en vit trappa.
En grupp män spelar instrument på en scen.
En kvinna på sin mobil, och en man som ligger bredvid henne på sin mobiltelefon också.
Folk i piratkläder spelar i ett band.
Ett barn bär hjälm rider en mountainbike mycket snabbt genom en skog.
Man på toppen av ett delvis fullbordat tak gör sig redo att lägga ner fler bältros.
En brun och svart hund vakar över en hört talas om djur.
En stor grupp poserar för ett foto på en gräsmatta.
Kvinnan går med sina barn och håller i glasstrutar.
Skateboarder i röd skjorta slipning längs kanten av en betong ramp.
Två tjejer spelar softball och en glider till hemmaplattan.
En grupp individer som chattar på en bar.
Byggarbetare balanserar på en smal bjälke långt över marken.
En pojke kastar löv i luften.
Svart, brun och vit hund hukar på tre ben i gräset.
Skateboardåkaren kommer upp på rampen.
Flera människor tittar som en skateboardåkare hoppar ner för en trappa.
En hund hoppar av en surfbräda
En pojke står mitt på vägen och sparkar en röd boll.
Ung flicka i rosa hatt tar bilder.
De leker med en fotboll på stranden.
Två män spelar i ett sportspel tillsammans.
En man i uniform bär hjälm med hakband och röd topp.
Den bruna och vita hunden går på grunt vatten.
En pugghund står upp på två ben och tittar över en stenmur.
En man cyklar i skogen.
En vit och brun hund leker i smutsen med en leksak.
Människor i Ghostbusters kläder står på en trottoar.
Kvinnor målar en stor rutnät målning av Afrika och andra delar av världen.
Två hundar leker i grunt vatten.
Tre vietnamesiska kvinnor paddlar sina båtar längs flodmarknaden på morgonen.
Ett par stövlar bärs av en kvinna med orange strumpbyxor.
En flotte paddlas genom en vitvattensälv.
En man och en kvinna som tittar över ett räcke.
Killar som dricker på en full pub, bara småpratar och tar en öl.
En kvinna som spelar minigolf och sätter upp en blå boll ur vattnet.
Ett litet barn i en blå jacka använder sin gula bleka för att vattna en växt.
En kvinna som hämtar bollar från ett minigolfhål.
En pojke med röd skjorta viftar armarna i luften när han tittar på en annan person.
En kille hoppar från stenar i vattnet.
Två små orangea och vita hundar är i snön.
En blå byggnad har rök strömmande ut medan en brandbil sitter framför den.
En person som bär en röd jacka håller i en öl medan en man i vit skjorta följer efter.
En kvinna med en svart och vit tröja som står på en gångväg.
En man i blå skjorta som cyklar genom en park.
En grupp människor klädda väl, utanför 2 bilar
Fem militärer i blå byxor med mässingsinstrument.
De övar för bandet för paraden.
Ett barn i hjälm spelar på en skateboard vid en lekplats.
En liten flicka blåser ut ljusen på tårtan.
En familj och en man i militärkläder tittar på en tårta.
Sex personer går upp för en blå ramp
En kvinna som rider på en häst i en hopptävling.
Två hundar springer på en strand.
En blond flicka har sin mun öppen, tittar bort från fotografen.
Två gamla killar sitter på parkbänken.
En hund springer genom ett gräsfält med gula blommor.
En man med solglasögon som går i en park.
Folk sitter vid bord bredvid häckar.
En grupp kvinnor får smink applicerat.
En kvinna i vit klänning sitter medan en annan kvinna blåser torkar håret.
Pojkar kastar en fotboll på stranden.
En man sover på gräset och täckt med en rosa filt.
En pojke med blå skjorta står framför gårdens utrustning.
En naken flicka täckt av målade blommor design rider en cykel.
Ett par klädda i formella kläder kysser vid en sjö.
En grupp människor står utanför nära ett grönt tält.
Tre preppy män står runt ett formellt middagsbord utanför.
Två vita hundar plaskar runt i vita vågor.
En man som visar en bok på US Army Yongsan Library.
En kvinna som visar en barnbok som verkar vara upprörd över innehållet.
En dam som läser en storybok.
Två små barn dekorerar muffins med glasyr.
Kvinnor sitter runt ett rum och har en livlig konversation.
Kvinnan tränar sin hund att hoppa genom korgar med hjälp av träningsutrustning.
En man i en byggnad som spelar horn.
En svart hund simmar i en stor pool.
En äldre kvinna i en folkmassa som knuffar en rullstol.
En flicka med kort svart hår och en flicka med långt blont hår poserar medan skridskoåkning.
Kvinnan med röd rosett går förbi en cykel.
En flicka som ritade en bild med en dam som hjälpte henne att stå bakom henne.
Små valpar i badkar får duscha med handhållet duschhuvud
En fågel landar på stranden nära många andra fåglar.
En ung flicka står på sanden vid en strand.
En hund som hämtar en käpp i vattnet.
En tjej i röd skjorta svingar på magen.
Ett barn hoppar över ett hål i marken.
En hund biter en annan hunds nacke.
Ett barn som rider en röd och gul karusell medan hans fötter uppe i luften.
Den lilla flickan i baddräkt står nära sprinkler och skrik.
En vandrare poserar på en klippa högt i bergen.
En man och en kvinna sitter i små möbler.
En man som bär färgglada kläder och medaljonger på huvudet slår en trumma medan han står bredvid ett litet träd.
En mountain bikeer gör ett trick på en skogsstig.
En svart hund springer genom snön med något i munnen.
De två boxarna är kvinnor.
En kvinna med långt svart hår trycker ett vitt mönster på ett blått tygstycke.
Två indiska kvinnor tittar över tyg.
En brun häst är i en konstig pose medan galloping utanför.
En gammal man med beige hatt som spelar på sitt svarta dragspel.
En pojke är på väg att hoppa i vattnet.
Människor samlades längs vägkanten och höll flaggans färgade röda, gröna och vita.
En bicyklist som utför ett trick över en kraftigt graffitierad vägg.
Ung flicka som borstar en häst med en handhållen maneborste.
Två flickor sitter framför en staty.
Flygplanet böljande rök och ser ut som det kan krascha.
En skjortlös man lagar mat på en utegrill.
En man i en blå skjorta som städar fönster från en sele.
Skateboardare gör tricks på en trappa bredvid spegelbyggnader.
En pojke i en randig oxfordskjorta poäng.
En ung flicka dumpar konfetti på en kvinnas huvud när hon ler.
En man hoppar i luften mitt på en väg.
En liten pojke i blå skjorta och kaki shorts leker på en lekplats.
Två flickor är i en skolkorridor.
En person i en svart tank topp spelar franska horn med andra människor.
En ung flicka som håller två vandringsstavar står på en klippa i en bäck.
Balettklassföreställning med lärare i närheten som hjälper dem att minnas sina drag på scenen.
Två män som är uppklädda går längs gatan medan en annan man stirrar på dem.
En man som hoppar i luften och gör en split framför en vacker byggnad i bakgrunden.
Två små barn skyfflar snö utanför ett lägenhetskomplex.
Ung man med uppvänd hår poserar med ung man med solglasögon och kvinna med glasögon
En svart hund hoppar över ett hinder.
En luftburen cyklist hoppade från en graffititäckt ramp.
Tre män äter mat på en soffa.
En grupp människor som sitter i ett rosa rum med ljus.
En man som står på en stege och pratar med en annan man som hänger ut genom ett fönster.
En man och en kvinna på scenen framför en dans.
En person som åker skateboard på en skateboardpark.
Flera ungdomar rider på en stor gul fair ride
Flera äldre män sitter på en bänk i parken.
En ung flicka som gör ett mönster för att designa kläder.
En grupp människor är utanför och tar en källa.
Liten asiatisk flicka och pojke springer mot kameran i motsatt riktning mot de andra människorna.
En man håller i en mikrofon i vita byxor.
En man valpar framför en vit byggnad.
En svart man sjunger in i en mikrofon.
En ung flicka fiskar med några äldre människor, kanske hennes morföräldrar.
Den här personen gör ett trick på sin cykel.
En vuxen kvinna och en liten flicka sitter vid vattnet i skogen.
En man med väst och slips på att uppträda inför en publik.
En flicka som bär rosa hatt och grå byxor klättrar på ett kedjelänkstängsel.
En brun hund ligger på ryggen och slåss med en brun och vit hund.
Det finns en man som kastar en baseball och har en handske sin vänstra hand.
En asiatisk familj sätter sig ner för ett mellanmål
En pojke i röd skjorta fiskar med tre av sin vän på en bro.
En liten brun hund som föder upp några får
En ung flicka i rosa klänning med något i handen.
En dansare poserar i ett tomt rum.
En knubbig baby med orange hatt stänker i en ytlig kropp av vatten.
En man håller ett litet barns hand när de vadar i en grund flod.
En liten pojke spelar ett racing arkadspel.
En eklektisk grupp utför sin konsert, komplett med huva dräkter.
En man, som bär alla svarta kläder, springer nerför gatan när en bil kommer mot honom med sina strålkastare på.
Två honor hoppar av gungorna.
En bild av en gångväg formad av två rader av kolumner.
Folkmassorna står utanför nära en brandgrop.
Det finns en skara människor av män, kvinnor och barn.
En flicka sitter på en gungtur.
En man i vit uniform rider en motocross cykel nerför en skogsstig.
Personen går ner i vattnet.
Turister njuter av en traditionell båttur i lång paddelbåt.
En ung pojke sträcker sig efter och rör vid propellern i ett vintageplan.
En man och en kvinna som går nerför en trottoar, bord med paraply uppsatt i bakgrunden.
En kvinna hoppar på en brygga vid vattnet.
En tennisspelare försöker träffa bollen.
Två barn leker med dockor medan vuxna tittar på dem.
En person gör ett trick med en skateboard.
Mannen i den gröna skjortan tittar upp.
En grupp människor är ute på vattenfarkoster mitt i havet.
En festival där musik spelas och människor samlas.
Många människor sitter i baren med drinkar framför sig.
Handikappad kvinna som står framför en Tartuffe-affisch.
En ung man i gul skjorta flyger från sin surfbräda in i en våg.
Några par sitter på bönor bredvid en pool
En man använder sitt finger för att rita något på sanden bredvid ett barn.
En person som ristar en hök ur en trädstam med en motorsåg.
Mannen i de rutiga shortsen bygger en stor sandskulptur medan två andra män begravda i sand tittar på under ett blått paraply.
En ung kvinna som utför en traditionell dans.
En liten flicka leker i en boll grop medan hennes familj tittar på.
En kvinna som borstar håret i badrummet.
En flicka som tar en bild med sin mobiltelefon av en stor grupp människor.
Folk kliver på och av och orange buss.
En mor och barn beundrar en enorm mjuk figur av en gris.
En kille i rött på en cykel i luften.
En vältränad kvinna i röda löparkalsonger börjar springa på ett spår.
En man i blå skjorta på en restaurang.
Folk går på gatan där en barrikad har satts upp.
Grabben gör tricks på en skateboard
En man ser ett barn gå nerför gatan bredvid järnvägsspåren.
Medlemmar av ett marschband och dansare i gul-fringade kläder uppträder på en idrottsplan.
En bandmedlem i svart, vit och röd uniform håller sitt silverhorn.
En ung man som parasailerar i luften över havet
En äldre man som går på gatan och tittar på varor.
En ung flicka i rosa klänning dansar när en kvinna blåser bubblor.
En person i gul hjälm på en blå motorcykel gör tricks.
En gata med många leverantörer som säljer produkter inklusive melon.
En kvinna väntar på ett tåg på en tom tågstation.
En grupp unga vuxna duschar utomhus.
Mannen ligger på fältet och läser en bok.
Två personer står framför ett vattenfall.
Tre personer leker i ett snöigt landskap, en håller en stor snöboll redo att släppa den på de andra.
En marschbandslinje står och väntar i full uniform.
En skara människor som surfar på en utomhusmarknad en solig dag.
Det är ett par som går genom en bondes marknad.
En liten flicka i rosa skjorta sparkar en blå boll.
Människor med svarta ballonger på dem klättra smuts backe
Två unga flickor är armbrottning i sitt hotellrum medan en annan flicka tittar.
En flicka hoppar på sängen.
Mannen med orange skjorta slipar på sten, han bär inte skor.
En indisk man som jobbar på en stenmur.
En hund står på stranden med en stor sten bakom sig.
Två barn som bär denim går på en landningsbana.
En ung kvinna klär sig flamboyantly för någon form av festival med mycket färg.
En polisman har en misstänkt som sitter på marken i hans förvar.
Tre flickor dansar i ett stort rum.
Två kvinnor deltar i en kampsport match.
Ungar hoppar sina cyklar från jordramper nära en strandpromenad.
En närbild av två kvinnor som står tillsammans.
En man i vit skjorta och slips pekar på en bild i en barnbok medan en liten flicka tittar.
Ett barn häller sirap på en snurrande anordning
Ett barn i en blomtryckt klänning är i ett fält av blommor.
En man i skateboard i en tom pool.
Kvinna med inte en massa kläder på att spela på telefon
En ung flicka på en lekplats drar i snöret på en rosa jojo.
En pojke som bär en transformers t-shirt står med händerna utsträckta.
En man och en kvinna kysser.
En kvinna cyklar på en stig genom ett fält.
En brun hund rullar i gräset.
Kvinnan som bär en svart och vit jacka och röda stövlar bär också hörlurar.
En grupp vänner som äter middag tillsammans.
Mannen står bredvid en gul byggnad med ett blått fönster.
En kvinna i en park med lila blus
En person som uppträder inför en stor publik som sitter på gräsmattan
Två flickor som ger en stor hund ett bad
En ung pojke som bär blå pyjamas och gula glasögon hoppar upp i luften.
Ett barn i blått med glasögon.
Två svarta bälten sparring, en sparkar den andra i ansiktet.
En diskjockey har en bild av Michael Jackson.
En stadsgata, utanför en klädaffär, med flera förbipasserande.
En ung pojke hoppar från en gunga.
En flicka med en pojke som står bakom henne kliver in i en simbassäng
Tre hundar springer genom en manikyrerad gräsmatta.
En kvinna arbetar i ett laboratorium och undersöker något i en petriskål under ett mikroskop.
En pojke på en skateboard i luften
Två kvinnor och barn äter glasstrutar på bron dekorerade med blommor.
Sparka upp sand, en beach volleyboll spelare hoppar för bollen.
En skäggig man på en mässa med svart tanktopp och rutig hatt.
En kvinna med mörkt hår bär en grön tröja.
Tre barn i vinterkläder med teleskop utomhus.
Connah Store där de säljer tobak, godis, tidningar och kaffe.
En äldre herre som har sitt högra öga diagnostiserat av en läkare.
En ung flicka med blont hår som håller i en rail
Kvinna sparkar huvudet av en annan kickboxer
Man bär pojkar kommer att göra pojkar skjorta vågor på kameran under gay stolthet parad
En hund hoppar och springer genom skogen och snötäckt mark.
Hunden simmar över vattnet.
En kvinna med långt mörkt hår tvättar disken längs en smutsig vattenpöl.
En Boston baseballspelare på slagträ
En flicka lutar sig mot en köksdisk och skrattar, med midjebandet på byxorna i grenen.
En muskulös svart man som dansar i korta shorts.
En gatuartist med gitarr spelar musik och begär tips.
Hästar med jockeys deltar i ett lopp.
En man i kostym och glasögon går på en trottoar.
Den unga damen går nerför gatan en vacker dag.
Två baseballspelare på ett fält, med fyra åskådare, och en publik.
Två valpar leker med en plastpåse.
Två små barn ler och ett pekar samtidigt som det håller något rött.
En kvinna som följer efter på en tennisträff.
En person är klädd i en svart väst och hatt med massor av blommor fästa.
En liten flicka rusar ut bakom ett träd.
En ung man i grå tröja tittar in i stan.
En brun fläckig hund går i grunt vatten.
En brud och hennes tärnor står utanför och tittar på en man som kommer klädd i mörk kostym.
En ung man med lila skjorta gör limbo i ett gymnasium.
En man klädd som en kvinna klädd i ansiktsfärg sitter bredvid en annan man.
De två barnen tittar på den lilla gula hunden på trädet.
En man håller en inköpskorg framför en skylt på fiskavdelningen som säger "Fishmonger"
Det finns en odlad anka och flera ankor.
En person simmar under vattnet i en pool.
En person i en kanot är forsränning i vilda vatten.
Två personer cyklar på en solig dag i ett skogsområde.
Det finns många människor utanför en stor byggnad.
En ung man med guld korta shorts och en svart topp går i en parad.
Folk vinkar från en buss täckt av regnbågsflaggor.
Ett barn som bär något i skjortan går i regnet på gatan.
En man klär ut sig på Hawaii vid en lokal parad.
En man utan skjorta står i en parad och bär ett blomsterhalsband av plast.
En man är skjortlös och täckt av röda märken.
En person med rosa hår och tatueringar på övre och nedre delen av ryggen.
Två gamla män som pratar på bänken.
En man som sitter i sand och håller i en liten staty av trä.
En mänsklig figur i en naturliknande dräkt som står i centrum för uppmärksamheten på en fest.
En kvinna i röd skjorta och flerfärgad hatt diskar i handfatet.
En hund blir besprutad av en slang.
En pojke i gul skjorta och blå jeans hoppar över träningspyloner medan två pojkar klädda i fotboll uniformer ser på.
Två flickor sitter utanför trappan och pratar.
En liten pojke i en röd t-shirt hoppar från en blå rutschkana på en lekplats.
Detta barn håller röda, vita och blå ballonger
En DJ snurrar skivor på en klubb full av folk.
Två barn springer förbi en dinosaurie i skogen.
Tre personer, två män och en kvinna, cyklar i en parad.
Flera uniformerade män som bär flaggor och vapen leder en paradkontingent längs en liten stadsgata.
En långhårig kvinna med solglasögon dansar med två andra personer i en parad.
En man i uniformsvågor och ler mot kameran
Folk är klädda i lila, blått, grönt, gult, orange och rött kostymer för en parad.
Sex personer spelar xylofoner i ett mörkt rum.
Ett konsertband visar patriotism och talang, genom klädsel, liksom deras musik.
Den här herrn uppträder sin "en man"-show.
En man i vit skjorta bär en trumma när han talar med två andra män.
En kvinna håller ut ett fredstecken under en parad.
Några personer med en flicka som står upp i mitten och bär en grön klänning
En grupp barn beundrar bilder som ligger i sanden.
En kvinna i ett vitt förband står vid en disk med skålar med mat och tittar in i ett annat rum.
En man hoppar över en vattenfontän.
En man och en liten flicka i en rosa livväst och röd flytapparat som simmar.
En man som leker med ett litet barn i en pool.
En man med glasögon och en grön skjorta sitter vid ett skrivbord.
En man dyker ner i en swimmingpool på hotellet.
En asiatisk kvinna springer på en stenig stig.
En kvinna närmar sig en klippas kant.
En man med gröna glasögon gör ett trick på sin skateboard.
En kvinnlig löpare i ett lopp
Killen med skjortan av har en del av Calvin Klein underkläder visar och han går bredvid killen i vit skjorta och svart kjol och svarta leggings.
En person som cyklar, gör ett mycket högt hopp.
Ett litet barn som leker på golvet med bokstäver gjorda av kviltat tyg.
En person som hoppar från en docka i vatten.
En kvinnlig polis står bredvid en kvinna klädd som Jokern i Batman.
Två personer går över ett snöfält.
Två människor slåss mot varandra i någon typ av karate, båda bär den typiska vita kläder med svarta bälten.
Bill Cunningham på gatorna i NYC.
En jonglör och en pojke i en topp hatt med ett svärd står framför en folkmassa.
En mörkhårig man och en liten pojke använder skruvmejslar för att arbeta på skärmdörren.
Ett barn som gör trick på en skateboard på en bro
En man deltar i en bmx ras.
Tre personer går förbi ett urval av varnande kottar på en trottoar.
Skäggig man i grå och röd skjorta drar ett rep.
En man klädd i vitt, inklusive shin vakter, gungar fladdermusen i en cricket spel.
En grupp på tre hundar går genom snön.
En grupp människor som hjälper varandra att ta ner en vit duk.
En man i vitt står framför en grillfest.
En flicka med brunt, lockigt hår använder en blå mobil enhet inne i ett rum.
En far och dotter kastar stenar i en liten bäck.
En man och en ung pojke är ute och tar en paus från att cykla.
Person som spelar piano som har sjöjungfrumålning på sidan
Ett flygplan flyger över berget och försöker släcka en brand.
Två personer släpar en gul flotte in i en flod.
En grupp människor i gröna skjortor skjuter en kanon i en parad.
En skateboardåkare utan skjorta tar sin bräda i luften.
En grupp på fem pojkar sitter på klippor nära ett vattenfall.
Unga vuxna samlas nära ett starkt ljus.
En ung flicka med kort hår väver på en vävstol.
En kvinna i orange skjorta väver.
En sidoshow skäller på en liten scen på trottoaren försöker ringa in kunder.
En blond kvinna med en röd ryggsäck i snön.
Två personer sitter på bänkar och tittar på varandra.
En man som rider på en röd cykel.
Människorna i vita och maroon kläder är i en träbyggnad.
En man i solglasögon använder en stor metallgrill.
En grupp barn viftar med en stor duk upp och ner.
Medan flera människor går bakom dem, ritar en man och en kvinna på trottoaren.
Två flickor kolliderar under ett snabbt tempo spel att fånga flaggan i en park.
Ett knubbigt, rödhårigt barn svänger ett slagträ mot en boll på en tee.
En man i röd skjorta går förbi en cykel.
Trummisen slår trummorna på en utomhuskonsert.
En kvinna med hatt leder en liten hund genom en hinderbana.
Två killar som spelar boll och gör ansikten.
En kvinna som får en styling klippt från en kvinnlig hårstylist.
Två liknande bruna hundar delar hålla en vit leksak medan de simmar.
En ung flicka i gul topp och en blommig kjol står på en filt och biter på en leksak.
Lilla flicka i gul skjorta, håller en vit hatt när hon sitter på en filt nära ett träd.
Hunden hoppar högt för gul boll när en annan hund väntar nedanför på gräs.
En man som kastar sig ner i vattnet där en dam väntar.
En bicyklist som bär en hellment rider nerför en brant ramp
Man med mörkt hår och skägg äter en knaprig mat objekt dricka kaffe.
En man som bär inline skridskor åker skridskor nerför en cementvägg
En pojke som gör ett ansikte medan han sitter i sin bilstol
Två tjejer sparkar varandra i kampsportsuniformer.
En man som håller i en väska och går nerför en lång trappa.
En grupp college studenter samlas för att spela Texas hålla em poker.
En man som hukar sig ner och försöker använda en maskin av något slag.
En liten brun hund springer genom snön.
En kvinna och två barn står framför växter.
Två barn och en man tittar på gräset bredvid en sjö.
En pojke har ett rött paraply på en lerig gård.
En ung man i blå skjorta går förbi en vit lastbil på en byggarbetsplats.
En man i jeans tittar i baksätet på sin lastbil för något.
En grupp människor ser på som en man pekar på en whiteboard.
En blond liten pojke står vid ett stängsel.
En man går in i en stor gul och blå varmluftsballong på marken.
Nära snöflingsskylten sitter människan medan en annan står klädd i bricka och hörlurar.
En person som åker vattenskidor i en flod med en stor vägg i bakgrunden.
En man med gitarr talar in i en mikrofon.
En folkmassa står på en övervattensbro med stadsbyggnader i bakgrunden.
En skallig, skjortlös man som klättrar.
En man står på ett tak torkdukar ovanpå flera cementhus.
Man och pojke bär flytväst i vatten poserar för en bild
En man tar en bild av en cyklist som utför ett trick i luften.
En fågel lyfter, omgiven av stora stenar
Två honor sitter och jobbar på en konstnärlig matta.
Ett barn sparkar ut luften på ett sportevenemang.
Den vita kranen söker efter mat i en damm.
En pojke poserar med en metallslev i varje hand.
Två barn i jackor som går nerför en grusväg och bär blommor.
En båt flyter i vattnet.
Tre personer drar ett rep på en bergssluttning.
Grupp av mödrar och unga kvinnor som går med sina barn.
En manlig tennisspelare hoppar i luften när han förbereder sig för att lämna tillbaka bollen.
En liten flicka cyklar på en grusstig.
En grupp barn på en trottoar med två klara kannor.
Mannen i rummet bär en morgonrock.
En man hoppar från ledstången i en utomhustrappa.
En kvinna med en färgglad halsduk går ut.
Två kvinnor som sitter på en träbänk längs en strandkant.
Person som gör en trick cykel flytta i en skatepark.
En dam som bär röda glasögon och en blommig skjorta talar till passagerare i en buss.
En pojke sticker ut en aligatordocka från ett bilfönster.
En man och en kvinna lutar sig tillbaka på en bänk utanför en butik.
En man går genom Brenmark Tools &amp; Fasteners.
En äldre man i grå skjorta står vid en byggnad som har kött hängande ut för att torka.
En familj sitter i en park medan fåglar flyger runt.
Hunden springer bredvid havets brusande vågor.
En man i cowboyhatt rider en häst runt en tunna.
Tre män arbetar utomhus i solen.
En kvinna i svart skjorta sjunger på scenen.
Män tävlar på en väg.
Två herrar i smoking spelar tangentbord och gitarr.
Ett barn och 2 år gamla som ligger på marken under en spelmobil.
En flicka med färgade randiga byxor som borstar tänderna bredvid en vit soffa.
I en UFC match, en fighter har den andra nere på duken och är på väg att slå honom med sin vänstra hand.
Nån som åker skoter hoppar på en wheelie.
En skallig man i blått rider en enhjuling på en asfalterad väg.
En musiker och en dam med brunt hår ska snart sjunga.
En man med ansiktsfärg på en clown håller en ukulele och munspel.
En man och kvinna skrattar medan de håller ett pris.
Mannen gör en kaströrelse, medan han står på stranden.
Två boxare slår varandra i ansiktet samtidigt.
En kvinna springer med en hund på ett gräsfält med träd i bakgrunden.
En grupp människor som reser i en liten träbåt.
Det finns en kvinna som håller ett barn, tillsammans med en man med en rädda barn väska.
En pojke sitter på en båt med två flaggor.
Ett litet barn som spelar TV-spel på en Nintendo DS.
En man i brun jacka håller upp ett gult föremål.
Mannen med excentriska kläder och hår poserar i en butik.
En grupp barn i turen som kallas "Frog Hopper".
En grupp av fyra vänner, som är skjortlösa, hoppar med glädje framför en pir.
En kille kör en go-cart på gatorna.
En man kastar en wheelie på en cykel på en stenig strand.
En man som sover i en stol på en trottoar i New York City.
En man som skateboardar på en skateboardpark som är täckt av graffiti.
Många sitter på en mexikansk restaurang.
Folk går genom en trädgård mitt i en stad.
En ung kvinna som sjunger och spelar gitarr i en föreställning.
En grupp människor rider kameler med röda sitstäcken längs en sandig strand, och tre personer är till fots.
En flicka i rosa rock kastar löv i luften.
En grupp på fem arbetare samlas runt buskar bredvid en McDonalds skylt.
En kvinna på en surfbräda rider en våg
Två män sitter på en bänk och tittar på en vattenfontän
En skateboardåkare i svarta kläder hoppar över en bänk.
En brygga över vatten med en palm i slutet och fem båtar, under skymning.
En svart hund hoppar över ett hinder.
En flicka och en kvinna går genom en gata och är på väg att passera en telefonkiosk.
En man spelar säckpipa.
En svart hund som hoppar i vatten i skogen.
Den här pojken, klädd i röd skjorta och blå shorts, springer.
En man i blå skjorta spelar ett unikt instrument som stänker vatten.
En kvinna lagar mat i ett hemkök.
En liten pojke med hatt och sandaler sitter på gräset.
En cyklist gör en volt i luften.
En liten pojke går ner en blå och röd glida och glida.
En ung flicka hoppar genom luften på en lekplats.
Två barn och en svart hund leker ute i snön.
Svart hund med röd krage stänk i vatten
En man i en blå t-shirt som sitter på en säng och stirrar på något underligt
Ett barn håller ett äpple i munnen
En man och en kvinna sitter, medan de arbetar på ratten i ett blått fordon.
En grupp afrikanska amerikanska flickor sitter tillsammans.
En enda röd lagspelare bryter igenom två svarta lagspelare, för att slå bollen
Damen söker sina restaurangers produkter på gatan.
En man som använder rullstol pratar på ett fält med ett par kvinnor.
En man som sitter vid ett bord arbetar på en dator.
En man i mörk hatt och glas sträcker sig in i en skål på ett bord fyllt med olika skålar.
En man som håller ett barn sitter på en sten utanför.
En man i orange hatt och orange skyddskläder är upphängd från en byggnad och städar en del av byggnaden.
En arbetare hänger i en hög byggnad med utsikt över trafiken nedanför.
En man med orange skjorta och hjälm är upphängd i luften.
Baby i ett bubbelbad, som hålls av en kvinna i en blå skjorta.
En man i orange hänger vid en kabel och gör lite arbete på en byggnad.
Två personer äter på en restaurang.
En man och en kvinna beundrar en ljusröd motorcykel parkerad utanför en restaurang
Ett ungt barn som cyklar på en kärrväg.
Två vuxna och två pojkar poserar med berg och en sjö i bakgrunden
En corgi går nerför en stig i en skog.
Köpare köper produkter från en upptagen livsmedelsbutik i Asien.
En flicka blir nerstänkt av en havsvåg.
En kvinna som står med ryggen mot betraktaren har en plyschleksak i huven.
En man som lär sitt barn hur man fixar kedjan på en cykel.
Två unga pojkar och en flicka bor hårt på en gräsmatta täckt med torra löv.
En hund trampar genom mörkt grönt vatten.
En man som hukar och sprejar målar ett öga och ett äpple som bär gummihandskar.
En massa människor i kamouflagebyxor springer.
Det finns unga män som spelar fotboll, en man har tacklats av en annan spelare.
Brun och vit hund hoppar över lila och vit bar.
En grupp människor samlades runt en väggmålning i ett urbant område
En butikstjänsteman väntar på några kunder.
En skäggig man och en flintskallig man som bär priser på en karneval.
En pojke i blå skjorta på en dator.
Svart hund nära en docka tittar in i grumligt vatten
En kvinna och en häst hoppar över en miniatyrbyggnad.
En kvinna i en blå tank topp äter en chili ost korv.
En man packar upp en kylare fylld med mat.
En kvinna i en blå tanktopp sitter vid ett bord.
En ung man som tittar på en pinne.
En ung flicka i en blå skjorta med blå jeansshorts griper tag i toppen av en vit stenblocksvägg.
En kvinna som sitter vid ett bord i svart skjorta.
En man med gul skjorta och svart hatt är på en stig i vildmarken.
En man hukar sig på trottoaren bredvid en liten flicka.
En liten pojke ler när han har ett blått paraply ovanför sig.
En kvinna reser med en stor bläckfiskskulptur på stranden.
Två honor står bredvid varandra och verkar vara oexciterade.
En flicka sitter på en klippa bredvid ett vattenfall.
Två barn med shorts klättrar upp på ett djungelgym.
En familj besöker en skog som turister.
En man med ryggsäck över axlarna går genom en skog.
En grupp människor som går på en stig.
En tatuerad man utan tröja arbetar på en ställning utanför ett fönster.
En pojke på ett däck med en röd hink på huvudet.
En vit fågel flyger från vattenytan.
Tre kvinnor som bär traditionella kläder gör de sista touchen på sina kläder.
Tre män i kostym står framför skyltar som säger Ford, Auto Alliance och Mazda.
En asiatisk man ler när han gör sig redo att slå en biljardboll.
En ung dam som bär en röd skjorta som rör sig i rullstolen.
Flera kvinnor dansar och hoppar runt.
En grupp människor njuter av att dansa i ett rum.
En tjej i rullstol med röd och vit skjorta har röda prickar över hela ansiktet.
En man som bär röd jacka och knähöga stövlar är flugfiske.
En mamma och dotter delar glass.
En person i grå jacka med en svart budbärare tillbaka tittar över den närliggande floden och bron.
Två barn svänger på en lekplats.
De rugbyspelare i rött brottas spelaren i gult till marken.
En man i svart skjorta sitter bredvid en kvinna som spelar gitarr.
En grupp människor står under en struktur, ler och dansar.
Ett förvrängt foto av en lekande hund på ett blomsterfält
En man åker skridskor nerför en trappa.
Flera rådjur hoppar ett staket in i ett öppet fält.
En person som bär hjälm börjar falla från en silverskoter.
Det finns en kvinna med en grön halsduk runt huvudet.
En man i röd skjorta tittar i bakfickan
Tre vuxna njuter av mat runt en grill.
Två män sitter ner och läser bredvid ett bord med mat på.
En grupp människor tittar på menyer i en vit restaurang.
Den vita pelikanen flyger över havet.
Skäggig vit man tar på sig en grön dräkt.
En ung person som dyker för att göra en fångst under ett spel av ultimata frisbee.
Någon är lila bär en skärm gjord av trä och mesh.
Kvinnor på stranden återvänder till sin bil efter lång dag
Pojke i luften på cykel
En skara människor står på en våt trottoar framför en byggnadsskylt.
En liten flicka i gul skjorta som bär en korg med blommor.
Två läkare hjälper en liten äldre dam i rullstol, medan en annan kvinna tittar.
En kvinna i blå skjorta pratar med en grupp barn.
Kvinnan i den svarta skjortan lämnar papper till barnen som omger henne.
En kvinna som står bredvid en tvättmaskin och håller en stor prickplåt.
En liten flicka i en blå hjälm klappar en häst.
En man gör sin bil redo för tävling.
Två män i vita skjortor som står under vad som verkar vara ett stort svart paraply.
En pappa och hans son leker med några legos i barnets sovrum.
En ung kvinna tar hand om personens fötter.
En äldre kvinna får blodtrycket kontrollerat.
Två kvinnor med armarna om varandra ler.
En kvinna och tre män poserar för ett foto
Flera lastbilar stannade utanför för någon typ av utomhusevenemang.
Två män sitter bakom en pickup.
En kvinna som bär koloniala kläder sitter på gräset och läser för en ung flicka.
En man servar en röd och vit varm stång dragster bil.
Race team i svart t-shirt service deras röda och vita bil.
En gammaldags bil kommer nerför gatan.
En man med en tatuering med en ärmlös kappa balanserar en enhjuling på hakan framför en byggnad.
En depåbesättning håller på att göra ett fordon redo för loppet.
En grupp män står runt en röd och vit rolig bil vid dragloppen.
Ett team står runt deras dragster.
En man i solglasögon sitter i en tävlingsbil med en utsatt motor.
Röd båt markerade GRAHAM tävlingar över vatten.
En racerbil kör iväg medan en man täcker öronen.
En fin röd och vit bil leds till på en kapplöpningsbana.
En vit man med svart hatt och blå skjorta sittande på ett staket och spelar gitarr
En indiangrupp ber på ett däck med vatten.
En kille som spelar fiol på gatan och fyra kvinnor lyssnar på honom.
En man med byxor spelar gitarr medan han är på scen.
En medelstor bild av en folkmassa som protesterade för att få hem trupperna.
En kvinna i bra form är pole-vacklande över en bar.
Två män lagar mat tillsammans med en metallskål, nära en hängande växt.
En man som ligger på gräset bredvid en liten sjö.
Greyhound hundar ras på banan, med # 8 leder vägen.
Mannen cyklar uppför tegelväggen.
En grupp unga pojkar i motståndarlag spelar fotboll.
Två unga pojkar i baddräkter promenad
En surfare som fångar en stor våg i havet.
En kvinna spelar fiol utomhus.
En liten brun och vit hund leker med sprinklern i gräset.
En ung fair-kinned pojke rider en lekhäst på en lekplats.
En grupp ungdomar njuter av en rättvis resa.
Flera gammalmodiga bilar parkeras tillsammans.
En man och en kvinna går förbi en röd bil med en silver huva prydnad
Folk sjunger med stora maroonböcker.
En solbränd och svart hund hoppar genom en vattenspridare på gården.
En massa människor på en show.
En stor grupp unga vuxna trängs in i ett område för underhållning.
Två personer klädda i karatekläder slåss.
Fem unga män på tre flottar flyter i en vattenförekomst.
Kiter fastsatta på hjulförsedda anordningar i ett fält
Det är många män som tävlar på sina cyklar.
Kvinna och man sitter bredvid sin gröna lastbil.
En baseballspelare undviker en boll med sitt slagträ högt i luften.
En svart hund som försöker para sig med en brun hund
En man med glasögon och en blazer står framför en skylt.
En kvinna som går på en trottoar och gör sig redo att korsa gatan.
En kvinna i vit skjorta står vid en Gwan Multipurpose Centre skylt.
En äldre kvinna gråter medan hon sitter i ett fönster.
En kvinna som bär en färgglad sjal på huvudet använder en symaskin.
Fyra hundar leker och hoppar i luften utanför.
Mannen i den färgstarka skjortan balanserar en kniv på armen.
En man som uppfostrar en ung pojke till en klarblå himmel.
Hörni, det kommer att bli en lång rad hemma så vi måste alla göra oss redo och jag menar oss alla.
En kvinna lägger ut papper på ett bord.
En man med långt hår spelar en akustisk gitarr.
En man står bredvid sin monter och väntar.
Mannen sitter ner medan han njuter av ölen.
Två kampsporter tävlar i en match.
En kvinna i svart klänning med solglasögon.
En man står på ena handen på en skateboardramp.
Två kvinnor står nära en dörr.
En vuxen och ett barn går förbi en modern byggnad.
En liten flicka tittar på en födelsedagstårta medan en man håller ett barn.
En asiatisk man grillar kött.
En asiatisk kvinna borstar tänderna framför en spegel.
En dykare poserar för kameran under vattnet och håller ett stort ljus.
En kvinna med blå hatt och blå skjorta med gul kjol målar en bild.
En cykelförare balanserar sin cykel på en räls.
En kvinna sitter och läser i en trädörr.
Någon i astronaututrustning är under vatten.
Den lilla flickan i den gula hatten är begravd upp till midjan i sanden på stranden.
En kvinna som skrattar som sin man har armen om sig.
En man i silverbil pratar på mobilen och en annan står på trottoaren.
Fyra personer står på en båt på sjön.
En man, kvinna och en annan man går genom ett gräsfält.
En man med blå skjorta håller ut armen mot en haj.
En liten flicka cyklar och skrattar.
En grupp människor går in på en idrottsstadion.
En kanna med röd skjorta och vita byxor står på högen.
En kanna står på högen.
Ledande sångare i bandet "Green Day", Billy Joe, sjunger en sång på scen med en ung pojke i bakgrunden.
Fyra personer står på en flotte och seglar iväg på vattnet.
En rad människor lämnar trottoaren och går in i en gul skolbuss.
Högst upp på läktaren och tittar ner på basebollarenan.
En man i röd mössa, gul skjorta och svarta shorts tittar ner på en stadion.
En underhållare gör ballongdjur för barn.
En kvinna som bär solglasögon lyssnar på en Walkman och röker en cigarett.
En kvinna och ett barn sitter i ett stort träd med stora grenar.
Ett litet barn som tittar på en kaktusträdgård.
Orange hund ser över axeln, nära poster på landsbygden.
En kvinna med röd halsduk, vit skjorta och solbrända shorts ger en ljudsignal till kameran framför bokhyllorna.
En man i hatt spelar entusiastiskt fiolen på en trottoar
Ett barn i en barnstol med en röd mössa som säger "kärlek".
En bild av en trottoar mellan en väg och byggnader.
En kvinna äter vid ett bord när folk går förbi.
Barn i praktfulla röda, vita och guldklädda dräkter som dansar i en parad.
Två små flickor, en på golvet, och en på översta våningssängen, visar upp sin prinsessa slott våningssäng.
3 mörkhyade hanar, två skjorta utan, är på ett gräsbevuxen område med träd utspridda runt omkring dem.
Folkmassorna samlades på en brygga med fartyget "evergreen" i bakgrunden.
En Tribe Warrior klädd med kulturkläder.
En ung pojke med mörkblå hatt sover på en bänk vid en terminal.
Stor kommersiell tegelbyggnad med byggnadsarbetare och tung utrustning.
En äldre man med långt vitt skägg och lerstövlar gräver upp lera för en trädgård.
En kvinna tävlar i ridsport ovanpå en vit häst.
En grupp barn som leker sätter svansen på åsnan vid ett relä.
En liten pojke på lägret, i en blå skjorta, kastar en fotboll.
En man utanför i kocktunika packar upp små gröna grönsaker.
Två män står i en elektrisk utomhuslift.
Fem män i svarta och gula kläder stirrar upp och en kvinna håller en cykel stående bakom dem.
En man står i en körsbärsplockare.
En man från en infödd afrikansk stam som tittar ut i fjärran.
Två män i gröna och svarta kläder rider högt i en korg kran.
En pojke med blå strumpor och röda byxor och en skjorta med fingeravtryck hoppar in i huset.
En man i svartgula karnevalfjädrar som spelar trummor.
Det finns två barn i badkläder som leker utanför bredvid några träd.
En man med baseballkeps åker skateboard.
Två män står på en klippa vid kanten av havet.
Byggarbetare är upptagna med att arbeta medan människor går förbi.
En flicka som bär en blå och rosa baddräkt kastar stenar i en sjö.
Kokar i en pizza salong kolla ugnen.
Mannen bär lila skjorta och svarta byxor, håller en kamera, står i en stads park.
En man med en drinkkopp pratar med en annan man.
Ett barn i en suddig skjorta som leker i en rabatt.
Ett barn ler och hänger på ett litet tåg.
En man i svart skjorta som bär ett litet barn.
En liten pojke sätter ett slagträ på pannan och snurrar runt.
Flera män och kvinnor sitter i stolar på någons bakgård uteplats.
Två tjejer dricker på en fest.
En man i svart skjorta och en kastad röker en cigarett.
En stor man på en fest, med en drink i sin högra hand.
En man ler för kameran med en öl i handen.
En man står nära en byggnad.
En liten flicka i rosa skjorta sitter vid bordet och dricker en milkshake
Två honor tränar på en strand.
Två vandrare vandrar över en sluttande bergssluttning med djup pensel i fläckar.
En pojke i grön skjorta ovanför något blått.
Två gamla skäggiga män rynkar av sig och tittar ut i fjärran.
En countrypublik på en festival.
Två poliser i solbränna står på sidan av en stadsgata.
Barnet i superman T-shirt skrattar.
En liten flicka i baddräkt medan hon äter en vattenmelon i vattnet.
Två kvinnor som har kul på en fest.
En man med vit hatt lastar grenar i en flishuggare.
En grupp vänner firar på en fest.
En kvinna i mörk skjorta håller upp en fotoklippning på en fest.
En man som håller i en öl ler med slutna ögon.
En man och en kvinna framför en spegel ler när han kysser hennes kind.
En berusad kvinna kramar en berusad man.
Två collegekillar poserar för en bild på en fest på kvällen.
En person arbetar på maskinen.
En ung person ställer upp i en basebollmatch.
Folk gick upp för trapporna med en enda fil.
En grupp åskådare tittar på en körföreställning.
De väntar i en trappa.
Man i svart smoking sjunger sin solodel i föreställningen.
En äldre kvinna i mångfärgade kläder som sitter bredvid en hög jordnötter.
En person utför ett trick i luften med en smutscykel.
En blond kvinna och en man i jeans sitter på en bänk utanför.
En person går upp för en vit sandig kulle mot den blå himlen.
Många unga människor sitter och lägger sig på filtar på ett fält.
En brun fluffig hund ligger i snön med sin gröna boll.
En grupp män spelar hockey.
En kvinna i brun skjorta knäböjer på gatan.
Lillgrabben tar nåt från en docka.
Barn leker i vatten och tittar på en jättebild av en persons ansikte.
En mans himmel på snö med berg i bakgrunden.
En kvinna i rosa tröja sjunger för en man i kostym.
En man med hörlurar står framför en affisch.
En flicka med flerfärgade ballonger står utanför mitt i en folkmassa.
En grupp färgglada kajaker paddlar genom vattnet
Ett blont, manligt barn som hoppar i luften på en veranda i trädgården.
En man i röd skjorta böjer sig över utanför en tom byggnad.
Tre tjejer som gör backflips på stranden.
En blondhårig bebis som sitter i sin stol och får mat.
En man med en öppen skjorta och glasögon som håller en mikrofon och en annan man i en bowlingmössa och rutig kostym med en rosett på ett instrument.
Ett litet barn som bär många ballonger.
En ung pojke njuter av att surfa när solen ligger lågt vid horisonten.
En man som klättrar på en klippa.
Två personer med cyklar stoppas för att försöka fixa kedjan på en av cyklarna.
En grupp människor i ett litet torg.
Ett litet barn undersöker tvålsuddar i händerna medan han tar ett bad.
En byggnadsarbetare skapar ett moln av damm när han arbetar.
En kvinna med brunt hår sätter rött lack på tånageln.
En grupp människor utför en pjäs.
Framsidan av ett mycket litet matställe på natten
En ung pojke matar en hjort med selleri bakom ett stängsel.
2 kvinnor sitter framför sina bord och säljer fisk på stranden vid havet.
En far och son ser en man svetsa på en staty.
Man sitter på en stol på fälten och snider en stadga som stöds av en trädstam.
En liten pojke leker på en lekplats med gungleksak.
Flera män i silverdräkter cyklar tvärs över en gata.
En afrikansk kvinna som håller ett barn i ett fält.
En kvinnlig servitör balanserar en bricka med en hand.
En lockigt hårig flicka fängslad av en fjäril.
En flicka med rosa hår och neonfärgade kläder svänger runt en rosa hulahoop.
En grupp människor är på en anläggning.
En man ligger bakom en vagn och försöker sälja olika matvaror.
Det finns en kvinna som kastar dolkar på ett mål, vilket är en morot.
Två män och en kvinna tittar på bilder i en tatueringssalong.
En kvinna i gult och svart klädesplagg åker skidor.
En uniformerad man lutade sig ut från en sidopilots fönster av ett stort amerikanskt flygplan för att tvätta cockpitfönstret.
Två atletiska män och två atletiska kvinnor springer genom en park.
Ett foto av åskådare som tittar på bandmedlemmar uppträder på fiolen.
Två kvinnor svänger på en åktur.
En grupp kvinnor lyssnar på en presentation av en kvinna i en labbrock.
Två personer sopar en grusmark.
En grupp kvinnor i långa, vita kjolar knyter näsdukar till huvudet.
Ett litet barn i bara underkläder dammsuger.
En brunettkvinna, som bär en brun långärmad skjorta, rodnar på kindbenen.
En grupp människor som dricker och pratar
Två män rabblar en byggnad framför en stor grupp människor.
Barn fyller vattenkanoner från en hink nära en swing-set.
Fyra kvinnor klädda i vita Midriff visar kläder flaxa en vit lakan i luften.
Två dansare sitter på scen med dramatisk belysning.
Pojken i svart och röd baddräkt hoppar ner i vattnet.
Fem barn går på en sandstrand.
Ett litet barn i grått och orange blinkar med ögat medan det håller i sig silverbestick.
En svart man som bär glasögon ristar en stenskulptur.
En ung pojke som plaskar i en liten uppblåsbar pool med en grön rutschkana bakom sig.
Lille pojke i en lekplats sitter på gunga set
En kvinna i en svart baddräkt som hoppar ner i grönt vatten.
En pojke i slutet av en glida och glida.
En man som bär blå overaller och en blå hatt, rider en liten hus dragen vagn.
Ett litet barn gungar på en stolpe på en lekplats.
Två gamla män spelar instrument, en spelar fiol och en dragspel.
Frukt och grönsaker står fint arrangerat med två män i ryggen.
En grupp människor samlas framför en biljettförsäljare.
Två flickor går, båda med en vit skjorta och blå shorts på.
Liten flicka som leker i en sandhög med bilar och människor i bakgrunden.
En skäggig man som bär en bandanna med skallar på håller i en kamera.
En liten flicka på ett bröllop har en bukett med apelsinblommor.
2 barn som hålls av en mor i en massa människor
Två kvinnor bakom ett nät på sina mobiler med två män sittande på en betongplatta på motsatt sida av nätet.
En ung flicka har blommor i ena handen och en korg med en båge i en annan.
Två pojkar gör tricks på sina skateboards på en skateboard park.
Byggarbetare passerar varandra på trottoaren.
De två männen spelar schack i parken.
Tre män och två svarta hundar.
Två byggnadsarbetare som bär orange hårda hattar står på platsen för motorvägen.
Tonårsdansare uppträder på en tävling.
En liten flicka i en grön baddräkt blir stänkt i en vattenfontän.
Någon form av firande förmodligen i en afrikansk stad.
Detta är tidsfördröjning fotografi med en person som rör sig ljus runt i ett mönster i mörkret
Tre män och en kollar hans mobil.
Ett band i vita hattar och handskar spelar med en stadion ett folk i bakom dem.
Två män uppträder orubbligt kampsport i en trädgård.
En man i en tung svart rock bär en tidning förbi en annons för en espresso.
En man tittar ner från balkongen från en stenbyggnad.
Unga pojkar klädda som sammanflätade soldater som går i en parad i regnet.
Folk går runt på en fullsatt plats.
En ung flicka går på vägen, medan hon bär en röd och vit klänning och skor.
Tre personer klädda i gröna fjäderdräkter dansar i en festlig parad.
En äldre herre säljer produkter ur bakvagnen som en kvinna tittar på hans produkter.
Två män i kostym, en sittande och en stående, har en diskussion medan de väntar på kollektivtrafiken.
Fyra tonåringar sitter på en bänk på natten.
En grupp män njuter av en fiskedag.
Grupp av är samlade i ett rum, de står bredvid en vägg.
En ung man hoppar sin cykel i en skatepark.
En flicka i lila klänning sitter på möbler med röda kuddar, medan leende för kameran.
En man bär en kvinna över axlarna på stranden.
Två killar sätter upp ett slags tak nära vattenbrynet.
En man med kamouflageshorts som justerar myggnät.
En man med skägg som står i vattnet bredvid en träplattform.
En kvinna med hatt läser sin bok.
Två män sitter på en pontonbåt och håller åror och bär hattar.
En kvinna i en solhatt ligger på ett stort svart rör.
En kvinna i en orange bikini övredel masserar en mans rygg.
Man i flyt i vattnet.
En man njuter av solen och den fria luften medan han seglar på en båt.
En man som bär en grön skjortskateboard på en gata.
En man ler när han sitter i ett badkar i ett badrum.
En man knäböjer vid en maskin.
En vit man med en öl sittande på en svart ballong i en park.
En man i svart hatt som knäböjer för att hugga en träbit.
En dam i hatt står bredvid en bil med soffa och innerrör på toppen.
En kvinna sitter på en soffa och läser en bok.
En grupp pojkar njuter av en dag vid bäcken.
I den varma solen har en oländig men välklädd man somnat.
Människan drar vad som verkar vara en trätavla med en matta på toppen av en ytlig vattenförekomst.
En kvinna i vit skjorta och svarta bottnar.
En MMA fighter slår ner den andra i mattan under en match.
Två män slåss i en MMA match.
Det lyckliga nygifta paret tar en stund att skratta och fira innan de skär sin bröllopstårta.
Unga människor som står och ler.
Två unga kvinnor i färgglada kostymer visar upp sina hulahoop färdigheter på en vänlig tävling under en lokal festival.
Två män spelar en lek medan andra tittar.
Två personer, en med rutig skjorta, och en med en vanlig ljusfärgad skjorta, springer på en balkong.
En stor orange buss stannar på gatan.
En man som bär avklippta jeans och gröna gympaskor sitter med ett ben korsat över det andra.
En man som sover på en soffa framför ett glasbord.
En man håller en kvinna i luften medan han är ute i bergen framför en hängglidare.
En man som går framför en orange och grön bakgrund.
En man tar tag i en stege medan hans fötter flyger i luften.
Tre personer slappnar av på en sjös kant som sitter nedanför snötäckta bergstoppar.
En magdansös med röd och guldfärgad dräkt står med armarna ovanför huvudet.
En man klädd i en röd och svart morgonrock sittandes på en dykbräda.
En man exploderar ur det mörkblå vattnet och sprutar vatten upp i luften.
Ett barn som står bredvid en väg med bilar som passerar förbi.
Tre hundar leker i snön.
Tre hundar leker i snön, med en stad i bakgrunden.
En man klädd som en clown försöker tvinga en lång ballong i en form.
Två arbetare i orangea skjortor tömmer en sopcontainer.
Många människor tar bilder med kameror.
Kvinna i rött skift och långa vita strumpor knäböjer på tennisbana.
Två unga män i ovanliga kläder hoppar i ett gym.
En massa människor som sitter utanför en byggnad på natten.
En ung flicka står framför en vattensamling med händerna ovanför huvudet och ler.
En ung flicka som bär hatt och halsduk klättrar upp för en pjäs i trä.
Tre män i stridsuniform sitter på tegelstenar med ett träd i bakgrunden.
En gul hund som springer längs en skogsstig.
Fem män i asiatisk inspirerade klädesplagg sveper om sina huvuden medan människor samtalar i bakgrunden.
En kvinna på en strand bär upp ett litet barn i vattnet
En kvinna med rosa bikini som dyker ner i en pool.
En flicka glider in i en liten vattenpöl.
En upptäcktsresande hoppar av glädje nära sin snöcykel vid kanten av en stor vattenförekomst i ett område täckt av snö.
En kväll pratade tre unga damer på gatan.
En pojke som sitter i dörren till ett hus i en slum.
Hunden hoppar över stocken med en käpp i munnen.
Två personer i hårda hattar och skyddsvästar som arbetar med kabel i ett gräsbevuxen område.
Arbetare installerar nya vattenledningar.
En kvinna i svart klänning står ensam och ser ut över en stad.
En dam som skär velveetaost och gör ett lustigt ansikte.
En ung pojke och flicka gömmer sig i högt gräs.
En blond kvinna med solglasögon på huvudet.
En mamma som håller upp ett spädbarn mot axeln i ett kök.
En äldre pojke som håller i öronen på en yngre pojke.
En barnflicka tittar på sina grannars barn efter en lång varm dag i Las Vegas i Nevada.
Kvinnan i grått håller en liten flicka klädd i rosa.
En asiatisk man med huvudet böjt sig i bön framför en gyllene staty.
Mannen i den gröna skjortan ler och håller i en yxa.
En man sitter framför en dator och tittar på papper.
En skjortlös man rider sin cykel, som sitter på framhjulet.
Pojken i grått ligger i snön medan han tar en paus.
Två män jobbar på en tegelvägg.
Det finns en stadion full av röda platser, en hejarklacksledare håller upp en skylt som säger ROCKS.
En idrottsman i gymnastiksalen gör sig redo att börja sitt gymnasium.
En ung, rödhårig pojke är klädd i en banduniform och spelar sitt instrument framför bandet.
Svart och solbränd liten hund som går med spetsade öron.
Fem ungdomar hoppar i glädje vid kanten av det tropiska havet.
En ung flicka använder en mopp och hink på golvet.
Två kvinnor undersöker ormbunksblad nära en bokhylla.
En man i arbetskläderna drar i snöret med lastbilen i bakgrunden.
En man i ett verktygsbälte styr en byggarbetsplats där ett stort föremål lyfts.
En man som spelar gitarr och sjunger.
En märkligt klädd man med en rutig kjol och knähöga svarta stövlar står mitt i ett trångt område.
En äldre man pratar med två andra män i en folksamling utanför.
En mörkhårig tjej som står framför ett band.
En man och två barn går
En man i röd skjorta som talar från en predikstol med en Mac.
En ung man som skateboardar på en räls.
En kvinna står på ett podi med ett bildspel bakom sig.
En man som undervisar om folsyra
En liten flicka med blont hår bär en klänning och en hatt som säger "Birthday Princess".
Fyra fartåkare tävlar på en isbana med spandexdräkter och hjälmar.
Fyra åkare tävlar i en snabbåkningstävling, och slår på banan.
En kvinnlig talare talar om GlamWiki.
En del människor och en hästdragen vagn står framför en restaurang.
Två personer går på en stig genom skogen.
En naken bebis som ligger ner med slutna ögon.
En ung flicka sitter vid ett bord och skriver.
En man klädd i hatt och blå rock rider sin cykel förbi en utomhus gao qui stand på en solig dag.
Ett barn använder en pekskärmsdator i en butik.
En dam tittar på en affisch med ett ansikte och flera skedar.
Kvinnor kollar in Ron Negros hårmaskot.
Folk testar en speldemo på en mässa.
Mannen bär röd skjorta och jeans på en atm
Tre bruksarbetare i orange uniformer och vita hjälmar arbetar nära en stolpe, med två av arbetarna är marken och en klättrar på stolpen.
En stor grupp människor sitter vid borden.
En man i en olivskjorta sms på sin telefon när han sitter vid ett bord i ett café.
En man med röd väst och svart fluga talar in i en mikrofon.
En äldre gent visar sin expertis i konsert på sågen.
Två munkar går tillsammans och funderar på livet.
Den här mannen tittar på en målning, med en pensel i handen.
En man med en stor röd skål går mot en brun åsna.
En man med skägg håller i en gitarr när han sitter framför en mikrofon.
En musiker spelar musik nära ett träd.
En man sitter på en pall, spelar gitarr och sjunger in i en mikrofon bredvid en fontän.
En pojke i grå skjorta med två överdimensionerade gurkor.
Blommor är bakom den fluffiga hunden som kommer upp för trappan.
En kvinna med lavendelskjorta bär en stor bunt trä.
En hund med brindlefärgad rock springer över gården.
En grupp människor sitter tillsammans vid ett picknickbord.
Det finns en unge i en blå skjorta och shorts med en hund.
En person som spelar på en repsving.
Här är en bild av en ung pojke som spelar i en golfortsby.
En man som bär en kortärmad skjorta hukar sig bakom en gul solros.
Många människor samlas runt ett högt träd som har en stege som lutar sig mot det.
Pojke klätterträd med alla säkerhetsanordningar fastsatta.
En man som går nerför en gata kantad av palmer.
Flera studenter tittar på en lärare i konstklass.
En kvinna dyker med sina första armar över huvudet när en annan kvinna simmar iväg.
Två män håller röda mikrofoner och vita handdukar.
De fyra människorna går i regnet.
Två kvinnor och en grupp män i grå skjortor på en klubb.
En vit skjorta med design av en dam kan ses hängande på en fullsatt marknad
Män och kvinnor som går på trottoaren utanför en marknadsplats.
En man med verktyg i båda händerna fokuserar på sitt arbete.
En mamma som sitter på en kullerstensgata och ger sitt barn en drink.
En grupp människor handlar frukt på en marknad för stadsjordbrukare.
En vit tältad fruktställ med flera personer som shoppar i den.
En glad ung flicka med brun tröja, rosa skjorta och blå jeans hoppar från en trottoar.
Flera män sitter vid ett bord med öl.
En kvinna som bär en blå tank topp håller en boll och tittar upp uppmärksamt.
En kvinna som står framför en docka med kylare.
En livlig motorvägsscen med en kvinna som korsar en korsning till vänster
Man framför en stor glasbyggnad.
En ung pojke spänner fast en mans ansikte framför en vattensamling som omsluts av betong.
En kvinna håller ett gråtande barn klädd i rosa.
En kirurg arbetar på en patient med hjälp av kirurgiska verktyg.
En kvinna sträcker sig utanför en byggnad som heter Vira Virou.
En indisk kvinna sitter i ett litet rum och designar vackra bilder på tyg för att göra filtar och liknande på tyget.
Två barn studsar på en studsmatta utomhus.
En man klädd i svart svepande bruna kakelgolv utanför en kakelaffär.
Fotbollsspelare sträcker sig som förberedelse för ett spel.
En fotbollsmatch spelas på en stadion fylld med åskådare.
Gatumusiker uppträder framför bänkar.
En huvud i en vit skjorta och bruna byxor står framför en monter som säljer olika varor.
Två personer är på sidan av en glasbyggnad.
En kille med blont hår står på en scen och spelar en röd gitarr med trummisen i bakgrunden.
En mörkhårig man som sitter vid ett bord med en bok och drinkar.
Brandmän släcker en stor brand.
En unge med en blå skjorta som klämmer tvål i handen.
En grupp äldre asiater samlas och spelar instrument i en park.
En man och två små barn slappnar av på en campingplats, äter framför en brand.
Ett barn stirrar ner över en grupp människor som är runt en brasa.
Stor brun hund tuggar på ben ligger ner.
Två pojkar i blå skjortor sitter på en bänk bredvid en skön åktur.
En gift man i kamouflage tittar genom ett gigantiskt metallteleskop.
Tre män i hårda hattar och solglasögon närmar sig en stor vit lastbil.
En man högst upp i byggnaden
En man med hård hatt pratar på en mobiltelefon.
Mannen som bär byggnadskläder sitter högt uppe på en byggnad.
En man i blå skjorta svetsar.
En man ger en annan ett föremål vid ett järnvägsbyte.
En gammal minivan målad för att se ut som Mystery Machine från Scooby-Doo kör förbi en vit byggnad.
En man är svettig efter att ha sjungit på scenen.
Flera unga män i en packad bil reser med däck bundna ovanpå sin blå bil.
Tre personer sitter runt en grill på hopfällbara metallstolar.
Två små vita hundar är på en gård och jagar en röd boll.
En röd suv med en kvinna inuti
3 personer i en bil med rallydekaler, utrustning på taket och en mongolisk flagga flyger.
En hane går sin hund nerför gatan.
En man, klädd i hjälm och blå jeans, föll av en tjur i leran.
Det här badkaret bor inte i det gamla huset.
Människor köper frukt från en monter som bär meloner, äpplen och andra frukter.
Passageraren håller i lasten ovanpå bilen.
Person i en röd skjorta står på gatan bredvid en bil med många dekaler på.
En man på en häst försöker att lasso en hund.
Tre personer sitter tillsammans på en soffa i ett hus medan två andra står på sidorna.
Tre unga män håller i trådarna
Man klädd i business casual klädsel spelar saxofon med resten av ett band.
En pojke i randig skjorta spelar trumpet.
Unga saxofonspelare väntar under en paus i en föreställning.
Två barn ler när de förbereder sig för att göra sitt stora plask.
En ung kvinna i vit skjorta och blå slips spelar trumpet.
Ett skolband av unga elever uppträder.
Tre flickor står framför ett musikstånd med trumpeter.
Två unga pojkar med saxofoner.
En kvinna med handväska går förbi en kinesisk affär av något slag.
Festivalbesökare har roligt med sina barn
Män och kvinnor gör yoga på stranden.
En skateboardåkare med röd hatt och grön skjorta som sitter på en skateboard och tittar på andra åkare.
En grupp jordbrukare arbetar tillsammans för att slutföra en växtrelaterad uppgift.
Fyra hundar på koppel går nerför en trottoar.
Två kvinnor uttrycker sina åsikter på ett politiskt rally
Två män i blå skjortor och sex kvinnor i balett.
En kvinna med blont hår går vilt nerför gatan.
Kvinnan bär bagage och dricker pratandes på mobilen.
Ett barn ger en kvinna en möjlighet att engagera sig i dess värld.
Två matarbetare som lagar mat i ett kommersiellt kök.
Ung kvinna i kort vit klänning som håller en korg går bland sanddyner eller hyddor.
En ung pojke som bär en stor klocka äter en glasstrut.
Bära ett hårnät och blått förkläde en kvinna förbereder sig för att kasta något i en cistern.
En blond bebis med en hästsvans rider en hink sving.
En tonåring i vit skjorta och flip-flops är i rörelse på gungan.
Två pojkar leker i vattnet.
Ung man med en blå skjorta på och rullskridskor utför ett trick från väggen.
Äldre pojke rullskridskor framför små barn på skotrar.
Sex buddhistiska pojkar går längs en väg i traditionella apelsinmunkar.
En man utan skjorta utför rullskridskor på en kurs.
En smaklös man som sitter på en stol med svart hatt läser en tidning medan han lyssnar på musik.
Två kvinnor ler mot kameran medan de njuter av sin lunch tillsammans.
Barn reciterar något från vitt papper.
Två barn tittar på antika lokomotiv i en utomhusmiljö.
En svart man som ligger på en bänk med huvudet på benet på en äldre herre som bär blå jeans.
En man med en kundvagn säljer varor på en livlig gata.
Två pojkar i svart står bredvid både en cykel och ett träd.
Tre personer ser ett vindband uppträda.
Två män i vita hattar och orange västar arbetar framför en byggnad.
En kvinna i en blå tanktopp som cyklar.
En man i blå skjorta och khakis spelar gitarr.
Fem män pratar i ett rum med datorer i.
En kvinna i blå jacka står och ler på gatan.
Flera uniformerade män spelar musikinstrument.
Två äldre människor dansar till musik i ett band.
Två kvinnor bär infödda amerikanska kläder bär väskor
Två asiatiska män sitter på trottoaren med sina varor bredvid dem.
En lama står vid sidan av gatan.
Ett berg som påverkades av de tidigare vulkanutbrotten i den sydvästra staden av ett hopp.
Människor färdas via åsna med sina tillhörigheter på ryggen.
Två kvinnor som sitter vid ett bord i en park ler mot varandra.
Två personer tittar över en dal.
En man med en vandrande käpp och en orange ryggsäck, går genom en dalgång.
Folk går på en grusväg.
En samling blå tält, varav ett står Exodus, är uppsatta i ett frodigt landskap.
En kvinna i en blå jacka knäböjer bakom en skål fylld med tvålvatten.
En kvinna ligger på trottoaren på sin campingplats.
En ensam vandrare med käpp som går nerför en stenig trappa i fjärran landsbygd.
2 män i vandringsredskap går nerför en stentrappa.
En vandrare tittar på bergen.
En vandrare går upp för en stig av stentrappor med hjälp av en käpp.
Två personer med ryggsäckar vandrar bredvid en hög grå stenvägg.
En kvinna med röd ryggsäck tittar på Machu Picchu.
En person med en grön hatt som ligger ner på marken.
En liten pojke leker med en gul bil på trottoaren.
En äldre människa på ett höfält.
Här är en bild på två män som går in och ut från en polisstation.
En man fiskar i havet.
Ett par dansar alfredosco klädd i turkosa toppar, damen hålls upp i luften med händerna sträckta uppåt.
En person som går framför en vit byggnad med blå dörrar och fönster.
Kvinnan bär en hatt som står vid ett bord vid en tegelgata mitt emot kameran.
En fotografs syn på en livlig gata.
Det grönklädda bandet spelar på torget framför kyrkan.
Två barn skakar hand i ett trångt område.
Folk sitter och en hund står nära en stor inhägnad i staty.
En kvinna syr linne.
En ung man som bär färggrann klädsel och hatt sitter i en hydda.
En kvinna som tittar ut mot en utsikt.
Två personer står bredvid en del förnödenheter i ett bergsområde.
En chaparral landskapsscen tom från människans bostad.
En kvinna i blå jacka och en blå hatt som dricker te ur en blå mugg.
En alpin entusiast tittar nerför en stig.
En dam med solglasögon som sitter på toppen av ett berg bredvid någon annan.
En person går över en stenad stig.
Den här mannen i röd hatt sitter på toppen av ett berg en solig dag.
En kvinna erbjuder bröd till ett par turister.
En dam som sitter vid sitt bord och försöker sälja sina varor på en öppen marknad.
En infödd kvinna som visar en dekorativ filt.
Ett litet barn flyger en gul drake med utsikt över havet.
En liten flicka ska till skolan.
Två barn, i färgglada kläder, leker på ett fält med en stor sten i mitten.
En man paddlar på en blå boogiebräda.
En grupp turister tittar på en uppsättning kolumnar ruiner.
En ung man övar tricks med sin skateboard på en cement trottoarkant.
En ung flicka i blå hatt och rutig skjorta står framför en stol som håller i en bakelse.
Folk köper och säljer färsk fisk vid stranden.
Två arbetare hjälper kunder på Sonoma Artisan Sourdough Baker-stället.
En man spelar ett tv-spel medan en annan tittar i bakgrunden.
En kvinna med ljusbrunt hår som spelar fiol.
Två personer lutar sig mot en stenvägg och tittar på landskapet.
En man som går i väg på avstånd längs en stor mur byggd av stora block.
Vandrare klättrar en stig i bergen.
Någon skär en tomat med en kniv på en skärbräda.
En man hjälper en kvinna med sin fiskespö bredvid en sjö.
En brun hund som bär nyckel leker i smutsen.
Ett överviktigt par klär sig mycket lättvindigt för att gifta sig utanför.
En överviktig man och en kvinna är utanför och lyssnar på en tunnare man som läser ur en bok en delvis molnig dag.
En man som sover på en vit plaststol på en trottoar.
En man svetsar något av metall nära många verktyg.
En man som ser en person dyka ner i en simbassäng.
En kille i shorts, en huva, och vänder floppar spelar inomhus putt putt golf och är för närvarande vid "penguin hål".
Några barn leker.
En kvinna som bär underligt färgade kläder checkar ut i en närbutik.
En hippie gör två cappuccinos.
Arbetare och traktor finns bakom betongbarrikader och bitar av trasig betong.
En man går förbi en byggnad på natten.
Tre personer i en pool gör ansikten på personen som tar deras bild.
Med fokuserade blickar stirrar tre unikt klädda skådespelare utanför scenen.
En kvinna bär på en ung pojke som håller i ett löv.
Cyklist som cyklar över en metallbro.
En man med hatt, vit skjorta och tröja knäböjer på en matta.
Två barn på gatan som tvättar sina ansikten.
En gammal man i rutig skjorta och blå byxor tittar i ett teleskop en solig dag.
En ung man hög i luften utför ett cykel stunt.
En liten flicka i en klargrön baddräkt leker i sanden med en blå spade.
Två personer med paket, gå på avstånd på en strand mot vattnet.
Två afroamerikanska män som gick förbi ett skyltfönster med en docka klädd i randig skjorta och randiga byxor.
Två kvinnor som beställde spannmål vid ett gatuskott.
En kvinna i brun rock och vit halsduk går på en trottoar.
Damen tar en bild i spegeln medan hon håller i sin utrustning.
En kvinna som håller ett äpple bredvid en uppvisning av apelsiner, äpplen och meloner.
Tre barn säkrar en segelbåt till en docka.
En man med vitt hår och ett vitt skägg i svart kostym tittar på ett papper i en kontorsbyggnad.
Omkring åtta kvinnor i lila och blå klänningar buga mot en man klädd i svart.
3 damer hoppar från en sten i öknen med berg som bakgrund.
Efter en sandstorm renade en underhållsarbetare skräp från de historiska ruinerna.
Två män och en kvinna står på stranden av en flod och kastar stenar.
En gammal man som står bakom en korg full av gröna stjälkar.
Två män är ovanpå en vit yta i en grumlig vattenfront inställning.
Kvinnan i en blå aftonklänning har en mikrofon på scenen.
En man med en vit klänningskjorta blandar kort bredvid en dam i en brun skjorta.
Två personer cyklar nerför en grusväg.
Två personer på en scooter väntar på att en man med gitarrväska ska korsa gatan.
En blond tjej i en gul och svart jersey spelar fotboll.
En brun hund bär ett föremål i munnen på en snöig bergssluttning.
Två män i vita och orangea overaller som hoppar fallskärm.
En kvinna i grön klänning som tittar på en annan kvinnas ring på en gata.
En pojke hoppar på stranden.
En grupp människor i en liten glänta av dött gräs.
En färgad pojke sparkar en boll medan två andra pojkar tittar.
En ung flicka har händerna i ett badkar med vatten med löv i.
En man i gul skjorta gör östasiatisk kalligrafi.
En hane går ut i regnet.
En ung man som bär lövverk på ryggen och klättrar i stentrappor.
Gammal man i tredje världen knäböjer medan han arbetar med en stor hammare.
En man som gör ett trick på en cykel medan han är i luften.
Tre kvinnor sitter på trappan och pratar.
En man som målar ett däck bredvid vattnet.
En man i vit rock står framför en marknad och kylare.
En man som sitter på en soffa klädd i blå skjorta och håller i en kamera
En stor grupp människor samlas runt två tåg på järnvägen.
En gammal man sitter på en terrass i solen.
Här är en bild på folk utanför som väntar på att den stora sjöbussen ska ta dem någonstans.
Folk tittar på när två tåg går på spår.
Två barn står på sina händer i en dörröppning, medan två vänner observerar dem.
Ung rödhårig, tittar genom ett guldfärgat teleskop.
En man i vit skjorta sitter vid en vit och blå dörr.
En man som sitter i ett rum med blå väggar under sömnaden.
En man med solglasögon, vit skjorta och jeans spelar minigolf.
Två barn leker på en strand, en i rosa, ritar i sanden och det andra barnet, i grönt, står i vattnet.
Två ungdomar går nerför en kulle på en rutschbana.
En kvinna går medan hon håller en liten pojke i handen.
En man och en kvinna äter en måltid utomhus.
Två kustbevakningsofficerare ute på ett träningsuppdrag.
En yngre pojke som försöker raka sig medan en äldre man i bakgrunden tittar på honom.
Två personer som bär vitt duellerar medan en publik tittar.
Ett hånfullt svärdslagsmål i något latinamerikanskt land.
Hunden bär en rosa tröja.
En rad män lutar sig mot en vägg som en man med ryggsäck går förbi.
Tre män arbetar under en het sol.
En man med svart hår har en gul penna bakom örat.
En person som håller en "Boombox" på toppen av en buss, eller båt.
En man i uniform håller en stor kamera vid havet.
En kvinna som leker med sin hund på stranden.
Ett stort antal människor står i kö på en snabbmatsrestaurang.
En man som cyklade uppför en telefonstolpe.
En man gör mekaniker på en sandbuggi.
De beväpnade SWAT-officerarna vaktar det avspärrade området medan de inspekterar en ryggsäck.
Tre personer med specialutrustning går över gatan nära en brottsplats.
Det finns folk som väntar på att checka ut i en affär.
Två män trampar på stenar för att korsa vatten.
Kvinnor i blå kjol framför ett träd
Polisen som rider i en stor taktisk för lastbil i ett urbant område.
En grupp människor samlas och poserar för en bild.
En blond-hårig läkare och hennes afrikanska amerikanska assistent såg ut att kasta nya medicinska manualer.
En kvinna som jobbar provar den nya gula jackan
En grupp kvinnor står tillsammans i en rad och tittar på böcker.
2 vita damer i casual kläder.
Fyra registrerade sjuksköterskor klädda i smocks peer ner i mobil bin fylld med diverse objekt.
Sjuksköterskor i en medicinsk miljö samtalar över en plastmugg.
Tre kvinnliga arbetare på en medicinsk anläggning som tittar på tryckt material.
Tre människor rider i en karneval twister rida.
En läkare och sjuksköterskor på ett sjukhus som står bakom en vagn
Två unga sjuksköterskor visar leksaker för barn att leka med.
Två sköterskor tittar på saker i en vagn.
Sjuksköterskor tittar på en bok om barn.
En blond kvinna i svart skjorta poserar med en gul stjärna och en bok.
En skara kvinnor står tillsammans.
En polis, och två kvinnor poserar för en bild bredvid en officerare fordon
En man röker en cigarett och håller i en honungskaka.
En kvinna i blå klänning och regnkängor moppar kullerstensgatan.
Någon som flyger med hjälp av en ljusröd och svart fallskärm.
En kvinna i svart och rött lyssnar på en Ipod, går nerför gatan
Livvakter som undervisar i simlektioner för lokala barn vid poolen.
En man i vit skjorta använder en svart tavla medan andra sitter vid ett bord och tittar.
Flera människor står på ett fält med utplacerade fallskärmar.
En man som ligger på marken med armen under en bil vit tittar på honom.
En man och en kvinna som går på en snöig stig.
En grupp barn och vuxna leker i en pool en solig dag.
En man som springer utan skor på fötterna.
En smal man som bär rullade byxor och en randig vit och blå skjorta går på sand.
En man säljer frukt på gatan från en vagn.
Det finns en grupp människor som står utanför en liten byggnad i en by
En grupp ljust klädda människor firar på en festival.
De två hundarna slåss ute i snön.
Pendeln läser tidningen när man rider på en båt.
En kille i svart skjorta ritar på en vägg
En äldre blond dam i vit skjorta korsar gatan.
En man som står bredvid en annan man och tar emot en check på 10.000 dollar
En skara människor står utanför bredvid en gata.
En kvinnlig lärare pekar ut något för en ung kvinnlig elev som sitter vid ett skolbord.
Två män, en håller en cigarett, sitter vid ett bord utomhus på gatan.
Två män klädda i en kamouflageuniform försöker fixa en motorcykel medan en tredje man står i bakgrunden.
En flotta av små fiskebåtar som kommer till stranden.
En ung pojke, som har blå skyddskläder på rullskridskor, är böjd över ett knä.
En man i svart hjälm som kör en röd ATV.
Olika frukter finns på en utomhusmarknad i vad som verkar vara Indien.
Två medelålders män med blå skjortor som pratar.
Två mosaikarbetare i vita jackor arbetar på ett noggrant utformat kakelgolv.
Tre personer står vid en röd kärra.
Bare bröst man med boll mössa sitter i en utomhus arbete butik
En massa män hjälper till att fånga fiskar.
En asiatisk flicka dricker en kopp kaffe i en restaurang bredvid ett gäng röda blommor i en gryta.
En smutscyklist rider genom en del sand som åskådare klocka.
Den bruna och vita hunden bär en mycket stor käpp över snön.
Två hundar i snön.
Han jobbar på en tekanna som sitter på golvet i garaget.
En man i en mauvedräktsjacka står nära ett fartygs hjul.
En fotbollsspelare följer motståndarna quarterback, som är på väg att kasta bollen.
En utsikt över en rak väg med en kvinna som joggar längs sidan.
Mannen i svart skjorta och Bugs Bunny slips visar konstigt ansikte med kondom över huvudet.
En kvinna som stirrar ut över ett räcke från en gångväg.
En hund som går längs sidan av ett hus i snön.
En man är midja djupt i en flod som kastar ett nät.
Mannen i den grå skjortan försöker laga en brödrost.
Folk går längs en sandstrand på en klar dag.
En leende ungdom i en blå skjorta poserar på några utomhustrappor.
En trottoarkonstnär som skapar sitt nyaste mästerverk med krita.
Ett par tupplurar i gräset framför parkerade bilar.
Man släpar en båt genom leran.
Flera människor handlar på vad som ser ut att vara någon form av gatumarknad med bilar och graffiti och gatukonst i bakgrunden.
Folk tittar på en gatuartist som gör tricks med eld.
En ung flicka i rosa skjorta som sitter på en docka och tittar på en vattenförekomst.
Två arbetare tar en vattenpaus.
En gammal kvinna i tyghatt syr tyg.
En brandman strängar nödsamtalsband.
En korthårig man med blå skjorta pratar med en grupp människor utanför pueblo huset som har en vit dörr och en balkong.
En man spelar gitarr på trottoaren nära en byggnad.
En man på en cykel är utanför en cykelaffär nära en rad cyklar.
Skyddsstoppning redo för någon typ av uppställning.
En gatubusker som bär en topphatt uppträder med eld framför en stor publik, en del sitter och en del står.
En man dricker en öl medan han samtalar med en kvinna.
En man håller ett blått fiskenät framför några stenar.
Tre tonåringar lastar av en lastbil med vattenmeloner.
En cyklist fokuserar på sin resa när han passerar en sjö omgiven av kullar.
Sitter i en strandstol och tittar på vattnet.
En man roddar framför en kanot i en stor vattenförekomst.
Två barn med blont hår leker på en blå bild.
En man i vit mössa målar en byggnad med sina vita markiser medan han tittar på den.
Man i vitt tittar ner läs med två män i bakgrunden.
Två män lutar sig ut genom ett fönster och tittar på något åt höger om dem.
En kvinna sitter bredvid potatis och grönsaker.
Ett ungt barn i blått sopar golven som sina föräldrar.
Två hundar leker med varandra.
En man i svarta byxor, vit skjorta som spelar flöjt som en dam i rosa danser
Man hoppar över andra män med en grupp åskådare.
En svart gruva rider en stor trehjuling med tre stora tunnor fastspända på baksidan.
Hunden jagar fåglarna ute på fältet.
En infödd kvinna är omgiven av korgar med färsk fisk som hon säljer på en lokal marknad.
Ett barn i en orange tröja håller upp en sandal och ler.
Ett barn står mitt i vattnet med armarna upplyfta över huvudet.
En trevlig omstridd fångst under en ultimat Frisbee spel.
Ett dansande par gör ett dopp där mannen hukar sig nästan till golvet.
En blond man i randig skjorta som pratar i telefon medan han kopplar av i en stol.
En kvinna i blå klänning sitter framför hinkar med hö och spannmål.
En man i blå skjorta och keps håller en liten afrikansk pojke.
Kameler stiger för att ta en passagerare från en vit sandstrand.
En grupp människor pratar utanför på natten.
En kvinna med blå topp och vita byxor som arbetar i en butik
En äldre kvinna håller i ett litet barn.
En kvinna som bärs av två poliser från en folkmassa.
En liten grupp män äter middag och pratar.
Sovande afroamerikansk kvinna som håller sin sovande son under en tågresa.
En person cyklar framför tegelbyggnader.
En man i allt blått som jobbar på ett tåg.
En liten pojke leker med några tåg.
En svart kvinna i vit skjorta och röda flip-flops håller en bläckfisk.
Två poliser väntar på tre äldre män.
En man som bär en vit skjorta och en hatt, rider sin cykel, gör en obscen gest till fotografen
En flicka som står på stranden håller upp en död bläckfisk.
Ett gäng dockor som sitter på ett bord med en liten flicka i en blå tröja som står bakom dem och ler.
Människor med promenadkäppar vandrar nära stranden.
Ett Mariachiband som uppträder på baksidan av en restaurang.
En man som badar sig i en fontän.
En äldre man i svart jacka och blå shorts sitter på en cykel.
Ett barn med vått hår håller en fjäril dekorerad strandboll.
Två kvinnor i identiska klänningar och skor med olika färgade hattar sitter på en bänk med en häck i bakgrunden.
Ett litet barn leker på en elektronisk enhet med en stilus
Barnen såg den unge pojken skriva på den orangea tidningen.
En server på ett matställe som städar bänkskivor.
Små barn kastar hö över ett stängsel mot en brun häst.
Konstnär i gathörn säljer sina konstverk.
En modedesigner arbetar på sin ena design i sin studio.
Människor som sitter på marken och tittar på en soluppgång eller solnedgång bakom ett berg.
Detta är en grupp kvinnor som tar hand om några korgar fyllda med föremål, möjligen frön.
Tre personer hoppar över en presenning, med en djungelbakgrund.
En man står ny en såg med en vit brevlåda i förgrunden.
Gruppen ungdomar befinner sig i ett bubbelbad och njuter av det.
En man leker utomhus med två hundar, varav en försöker fånga en boll i luften.
En kvinna cyklar mot rött ljus.
En äldre man som bär solskyddsrock cyklar nerför gatan.
En cykelcyklist med en blå ryggsäck som går över en bro.
En man som surfar på stora vågor med en klocka på.
En flicka i en vit tank topp rör sig för att någon ska komma närmare.
En man och en kvinna som kysser varandra på en tågstation.
En kvinna i pionjärklänning sitter vid ett bord.
Man i en färgstark sombrero och poncho sitter på gräset med 2 getter och en lama.
Två unga män sitter vid ett bord och ler.
Unga flicka läser beskrivningen av park staty; det finns träd i bakgrunden.
En grupp barn går nerför en rad håller ballonger.
En man som använder käpp går över de vita linjerna på en korsning.
En grupp män spelar schackpoolside.
En man tar ett foto av ett par som står bredvid en skulptur utanför.
Två bicyklister rider förbi ett brunt fält.
Två äldre pojkar och två yngre pojkar tittar ut över vattnet medan de är på en båt.
En man spelar dragspel på trottoaren framför en affär.
Två flickor som sitter i gräset och bär hatt äter snacks.
En äldre kvinna plockar upp mat ur en kastrull.
En kvinna i gul skjorta med ljust orange hår avdelar från en ölkran.
En surfare rider på inkommande vågor längs stranden.
Två män surfar på en liten våg med en stad i bakgrunden.
Barn och deras föräldrar klättrar upp i ett metalltorn.
En actionbild av en volleybollspelare som spikade bollen.
En man kör en blå motorcykel.
En ung flicka med en saknad sko hålls av en kvinna i vita byxor med en svart topp.
Ett blond barn som äter en muffins med blå glasyr.
Bilden är att fyra män spelar på ett utomhusbröllop.
En tennisspelare visar en tvåhänt förhandsskott under en match.
En surfare som bär våtdräkt och använder en ljusfärgad tavla fångar lite luft.
En kille i rutig skjorta som går med en svart väska hängande från axeln.
En man och en kvinna på en bondgård bakom två tjurar.
En liten pojke skyfflar snö.
En dam med glasögon och en blå skjorta med axelväska är på väg att ta en bild med sin kamera.
En man och en kvinna reparerar något.
En parasailer hänger på bogseringsrepet.
En vindsurfare surfar på skumma vågor.
En man och en kvinna, båda knuffar barnvagnar med barn i dem, stoppas och tittar på varandra.
En man som håller i blommor medan en hund sitter i en cykellåda.
En man är upphängd i luften på kablar medan han gör lite arbete på en byggnad.
En hund som springer med något i munnen
En man i blå skjorta sjunger medan en flicka i svart klänning spelar gitarr i bakgrunden.
En person står i kostym på en gata.
En man och kvinna förbereder en blandning framför en rad cyklar.
Pojke i röd skjorta klättrar upp för en blockvägg.
Flera israeler står mitt i en upptagen korsning.
Man klädd som Darth Vader spelar en fiol på trottoaren.
Sex flickor dansar i en rad på ett idrottsevenemang i ett gym.
Brun och vit hund med baseball i munnen.
Den här personen är på väg att sätta papper i en kopieringsmaskin
En man i röd skjorta spelar pool.
En grupp unga kvinnor som bär blå tank toppar och vita kjolar alla gör en synkroniserad jubel.
Barnet får mat på en sked
En flygvärdinna serverar gods till flygplanets passagerare.
Två män spelar scen när de är klädda i karaktärskläder.
En flintskallig målare som arbetar på en bit på gatan på dagen.
Två personer kysser varandra på en gul linbana.
En man håller ett barn inlindat i en handduk på axeln.
En äldre manlig frisör som rakar en annan mans ansikte.
En ung man i svart jacka och svart keps spelar trumpet.
Ett band repeterar i sitt garage.
Musiker står på scen med sina instrument när en rad människor står framför dem.
En man i en grön skjorta sjunger in i en mikrofon.
Tjej i röd och svart skjorta som sitter framför ett tangentbord och uppträder med andra bandmedlemmar.
Två tjejer pratar på en fest.
En man och en kvinna som står utanför ett hus bredvid en ljudhögtalare.
Flera personer håller behållare med alkohol i ett rum.
Unga vuxna konsumerar mat och dryck bredvid tvättmaskinen.
Två personer på en fest eller konsert
En man med guldhalsband, en röd jacka, ett örhänge och eyeliner röker två cigaretter samtidigt.
En man och en kvinna sitter på en bänk och spelar stränginstrument.
En glödande byst sitter mitt i ett runt bord med papper prydligt utlagda.
Tre bruksarbetare på en telefonstolpe.
En kvinna sticker ut huvudet ur sitt tält på sidan av en snöig moutnain.
Kvinnan klättrar upp i ett snötäckt berg och tittar på folk bakom henne.
Mannen bär en stor ryggsäck medan han vandrar genom snötäckt terräng.
En vandrare klättrar upp för ett snöigt berg.
En grupp människor trängs runt några trappor av en nöjespark.
En walmartarbetare som bär vit rock.
En man i en kontrollerad grön skjorta sitter ner och tittar på sina händer.
Några män sitter runt ett bord.
En brun och vit hund står på bakbenen och sträcker sig efter en boll.
Leverantörer i Europa, en man och en kvinna som förbereder sig för en dag med att sälja grönsaker och frukter.
En rödhårig dam och en brunettfärgad dam står nära en vattenfontän.
Mogna män med en gåva i knät medan ett litet barn öppnar en annan gåva.
Ett barn som sover som person har en bok.
En man Rollerblade över en gul stolpe på natten.
En kvinna står nära vattnet, ser ut att kasta något.
En man hänger på en häst när den hoppar runt.
En ung man på rodeoarenan bär cowboykläder på en häst som bär rep.
Ett barn med lekredskap är på äventyr utanför sitt hus.
En ung flicka i svart klänning håller en röd flagga och täcker ett glatt uttryck.
En man klädd i medeltida kläder sitter på en medeltida typ vagn.
Den lilla hunden hoppar i luften mot kvinnans hand.
Folk köper mat från en tillfällig matförsäljare.
Tre män sitter på en gångväg.
En man häller något från en burk på en smörgås.
En man och kvinna sitter vid ett bord i en restaurang med utsikt över bergen.
En kvinna sitter på en blå bänk och läser en bok.
En pojke med blå t-shirt, khaki shorts och sandaler går ut.
Man i blått och gult tittar på en Jumbotron.
Elever i en klass utför labbexperiment medan de bär glasögon.
En man i röd kappa som rider en vit häst i sand.
Upprörd kvinna i blå klänning som går i en stad.
En säkerhetsvakt står ensam vid en vägg.
Tre barn, som bär gröna, gula och blå uniformer, sitter och står nära två kvinnor.
En grupp barn, med vuxna hjälpare, arbetar tillsammans.
En ung pojke höjer handen, som andra unga barn skrattar i ryggen.
Tolv barn samlas på en utomhus tropisk plats.
En grupp unga asiatiska kvinnor som ler för kameran.
En kille som går uppför trappan och håller i en portfölj och en bok.
En person klädd i en röd huva sitter på en bänk med huvudet nedåt och lämnar över ansiktet.
Två barn sitter på trottoaren.
En ung man i vit skjorta håller båda händerna ovanför huvudet.
Två små flickor som läser och ett barn som lyssnar.
Åskådare klädda i ljusfärgade kläder tittar på när man klädd i vita byxor och barfota blåser en boll av eld.
Folk på en fullsatt tunnelbanebil.
Två stora bruna hundar springer genom snön.
Ett litet barn som leker med en volleyboll nära en vattensamling.
En man med en öl och hammare i händerna slår något på en rund plattform framför sig.
Fyra personer med hattar som sitter och äter på en bänk.
En liten pojke som ger en liten flicka en tröstande kram.
Två manliga brandmän med vita hjälmar stående framför en byggnad.
En man i vit kort och shorts träffar en tennisboll.
En tjej i vitt spelar tennis.
En kvinna i vit klänning och vita skor som spelar tennis.
Tjej i röd skjorta och vit tennis kjol lämnar tillbaka tennisbollen.
En kvinna, som bär flera mångfärgade hinkar tillsammans, sticker stenblock vid vattenbrynet.
En kvinna representerar University of Phoenix vid ett visningsbord.
En grupp människor rider på en rakettema nöjespark.
Pojke i grön hatt reagerar på historisk fläck.
Två anställda ser på som en annan anställd kastar deg i ett kommersiellt kök.
Pojke i randig t-shirt går längs en avsats.
Fem personer är jämnt fördelade längs ena sidan av en tråg full av ananas på ett stort fält.
En samling grönsaker sitter i korgar.
En mountain bikeer klädd i skyddande redskap rensar en liten smutshög på ett spår medan en publik tittar.
En ung kvinna sitter på en moped framför ett café.
En gatuförsäljare i en röd skjorta och vit hatt som säljer italienska Ices från sin vagn.
En man fixar en stege för att klättra upp och ner.
En man närmar sig en fallskärm som han kanske bara brukade landa på marken.
En kvinna som leker med en liten pojke på dragspel på ytterdörrens trappa.
Hunden bär en röd keps och har munnen vidöppen.
En knubbig man som går nerför trottoaren.
Tre män fiskar vid kanten av en betongbarriär som är byggd längs stranden.
En ballerina i svart klänning och tights dansar framför en betongvägg.
En japansk kvinna städar en byggnad från ett museum.
En cowboy visar upp sin mulåsna bredvid en häst som kör trailer.
En man i lila skjorta som spelar trummor framför en folkmassa.
Byggherren lägger upp stora betongtrappor.
Fyra män i tajta kläder, tre i blått och en i svart, justerar sina kläder medan de står på en asfalterad yta.
En man i jeans jobbar på ett gammalt tåg.
En orgelspelare sitter och leker inne i en kunglig kyrka.
En man i gul grävmaskin på en byggarbetsplats.
En liten grupp människor solar sig på spån vid sjön eller havsstranden.
Asiatiska Greyhound köpa resa någonstans.
En man och en kvinna läste i en kyrka.
En stor svart hund har tassen på en liten brun hund.
En man med hatt och hängslen går genom majsfält mot en silo i bakgrunden.
En skara människor utanför ett kinesiskt tempel.
Tre leende kvinnor klädda i svart följer en fjärde kvinna med tatueringar runt ett rep.
Två personer som använder en vattenbuffel för att odla ett vattnigt fält.
En man i blå jacka och rosa skjorta sjunger och spelar gitarr
En liten flicka bär rosa byxor.
Den stora, svarta, löparhunden har en rem runt bröstet.
En vit hona är ute på en marknad och tittar på frukt.
En ung pojke med ljusbrunt hår som sätter ansiktet i sin måltid.
En pojke i en grön och vit randig skjorta ser utmattad ut när han springer
Kvinnan i röd rock köper något från en gatuförsäljare.
Flera cyklar parkerade och ett par går tillsammans.
Tre män vid ett bord medan en tittar på att hålla sin martini.
En brandman som ska släcka en bilbrand.
Mannen i brun jacka med armen runt personen i svart jacka på blomsteraffären
Två personer sitter på en bar och pratar.
Åskådare tittar på, och en knäpper ett foto när en man hoppar från en bro.
En man som bär ficklampa på huvudet har handen i en rullväska med vajrar.
Tre tjejer spelar basket, nummer 35 håller i en orange, vit och svart basketboll.
Eleverna verkar vara i ett laboratorium.
Två killar, på i en maroontröja, den andra i en ljusblå, sitter skjortan och spelar tv-spel.
Två kampsporter med skyddskläder som slåss inne i ett gym.
En ung man blir flygfödd medan hans skateboard snurrar under honom.
En man förbereder sig för att sätta på en smörgås ombord annonsera en Ebay verksamhet.
En kvinna i en maroonskjorta förde samtal med en annan kvinna i en solbränd blazer.
Person i orange kläder liggande på en vägg
Grå och vit hund med röd sele och koppel går över en stenvägg.
En kvinna i lila skjorta bär tre fulla shoppingväskor.
En grupp människor går framför ett berg.
En man som bär en gul och svart hoppare gör akrobatik.
2 personer med ryggsäckar är vid ett bord med en kvinna med en beige blazer sitter bakom den.
Mannen i kostym sitter bredvid väggen av VHS tejpad.
En kvinna med glasögon sitter framför sin laptop i ett bibliotek.
Flygbolagskunder väntar på sitt bagage vid en bagagekarusell.
En man som rider en fyrhjuling genom leran och han ser väldigt lycklig ut.
Asiatisk kvinna håller flagga med kostym drake i bakgrunden
Två killar, en i gul skjorta och en i vit skjorta, leker med en Frisbee.
Svart kattunge äter en mal och ett blad.
En man i en röd tanktopp mediterar.
En kvinna med sandaler och en grå kundvagn som köper mat.
Bicyklisterna gör sig redo för loppet, greppar för sina cyklar, deras ultimata verktyg för att banka sin väg till mållinjen i detta lopp.
En ganska kvinnlig nyhetsreporter som filmas för en show.
En skara människor med parasoller står framför en röd byggnad.
En man utan tröja cyklar.
En man i jeans och en blå kontrollerad skjorta värmer metall med hjälp av smeds verktyg.
En asiatisk bicyklisk matförsäljare väntar vid korsningen.
En kvinna som bär en vit labbrock håller upp sin burk med en vit handske.
En man i blå skjorta jobbar på en cykel.
Mannen står upp och ner på flaskan, med händerna på marken.
En man som gör ballongdjur på en gata.
En grupp vandrare går en stig som leder från en sandstrand mot en kulle.
En medelålders man i kostym sitter på golvet mot en vägg medan han granskar sina anteckningar.
En byggnad som arbetar på en dimmig dag uppe i luften på en hiss.
En besättning gör någon redo för bungyhoppning.
En kvinna leder en oxe dragen vagn, med en man som går bredvid henne.
En kvinnlig soldat i glasögon visar ett föremål för barn.
En brunettkvinna i en blå satindräkt håller en slägga mitt i skogen.
En äldre man kastar plastpåsar nerför en trappa, attackeras till ett plan.
En gatumusiker som sitter och spelar gitarr med ett öppet fodral och en skylt som läser "Berätta varför MUSIC SUCKS".
Fyra elever poserar för en bild inne i ett klassrum.
Två personer är på gatan, och en har en cello medan en annan håller i ett dragspel.
Sveral ung man hoppar nerför gatan
En grupp människor som bär hattar och använder käppar går genom ett skogsområde på en stig.
Liten flicka spelar ovanpå en svart järn maskin.
Person på cykel håller en spade bredvid en kvinna i en grön skjorta med en tvättkorg på en dockvagn.
En mörkhårig kvinna tittar på en Apple laptop dator.
Två män i röd uniform och en blå uniformsstrid i karate i gymnastiksal.
En kvinna håller en liten pojke på en soffa.
En kvinna hoppar över en parkbänk medan hon kastar löv i luften.
En man som gör ett headstand framför orangea och vita barrikader.
Folk väntar på tunnelbanan på utomhusplattformen.
En brud och brudgummen går på en stig genom gräset medan ett annat par följer efter dem.
En man sparkar en bräda ur en annan mans hand.
Folk sitter i ett rum och pratar med en panel.
En grupp människor, av vilka minst två dricker ur vinglas, står i en korridor.
Tre ishockeyspelare i svart spel utanför.
En ung pojke klädd i vita shorts simmar under vattnet med slutna ögon.
En kvinna i grön skjorta håller i ansiktet.
Två vita kanopier med män som står under dem medan en man går sin väg.
En man fotograferar en bergsäng, med toppar i bakgrunden.
Två personer som bär uniformer och väskor går nerför gatan med en vägg i bakgrunden.
Två kvinnor sitter bakom sin monter på en gatumarknad.
En skara människor tycks lyssna till en talare medan en man och en kvinna talar bakom dem.
En mor och hennes två barn som knyter band över middagen.
En kvinna som bär glasögon och en svart blus håller en slev och en skål i händerna och klibbar en plastgaffel i tänderna medan hon står i ett kök.
En kvinna tittar in i en svalare glass.
En man med en kamera på halsen står utanför ett café.
En man i blå skjorta skär upp sin mat.
Två personer sitter på en bänk och njuter av naturen när ett stort moln tornar upp sig.
Skater sitter på botten av en skate skål med sin bräda.
En ung kvinna sitter på golvet och övar på arabiska bokstäver med hjälp av ett bläckhorn.
En grupp människor klädda upp för halloween.
En man med en ärtgrön jacka, vit hatt, solglasögon och en cigarr som går nerför gatan med andra människor runt omkring honom.
Kvinnor står bredvid ett produktionsstånd.
En man med vitt hår och ett långt vitt skägg äter.
En brun hund på koppel går i snön.
En enda hane som bär en långärmad vit skjorta som rider på en smutscykel.
En man i en blå skjorta som leker med rep i ett skogsområde.
En man i blå hatt och rutig skjorta stöter bort sidan av ett rockansikte.
Tre personer tittar på varor från en juvelkiosk.
En man med en grå jacka och vit hatt böjer sig över vattna en trädgård med en vattenbehållare.
Man ser sig omkring i ett konstgalleri.
En blå lastbil med lastsäckar på taket är på väg nerför en väg.
En kvinna som borstar tänderna.
En grupp på sex kaukasiska män står på byggnadsställningar och skrattar, dricker vatten och fotograferar.
Fem unga, stiliga män som hänger utanför byggnadsställningarna.
En ung flicka i en park undrar högt om vattnet vid fontänen är återvunnet vatten.
En äldre handikappad man sitter på en stol och håller i en flaska vatten.
En gammal man som läser en tidning på en restaurang.
Scubadykare undersöker ett havererat flygplan.
En trick ryttare bär en ljusgrön outfit som bär en amerikansk flagga ridande en målarhäst med grön ridutrustning.
Två mycket välklädda kvinnor står bredvid varandra.
En man i vit sjömansdräkt och flera andra människor drar i rep på ett segelfartyg.
En byggnadsarbetare står vid en stor lastbil och orange kottar.
En ung man i en lila amerikansk fotbollsuniform försöker anspela på en annan ung mans tackling i en vit uniform.
En man vilar på marken med en kopp.
En man flinar och håller upp en vit kaffekopp medan han sitter nära ett träd.
Fyra män pratar med en lastbil.
En liten flicka, som står vid sidan av vägen, tittar på en liten pojke medan han sitter på gatan.
Två män gör ett tillkännagivande på en balkong.
En tjej med en röd peruk ler som en massa människor klädda som clowner går förbi.
Två hundar leker på stranden tillsammans.
Klädda deltagare kastar konfetti och godis från en flotte under en parad.
En surfare som rider på en liten våg.
Två män står på en gata i en stad och mannen på rätt punkter på något.
En grupp ungdomar lägger händerna i luften i en livekonsert.
Mannen sträcker sig över bordet för att få mer mat.
En man som bär handske och slipar en bit metall.
En man med skägg spelar akustisk gitarr på gatan.
En äldre man sitter på ett café och kopplar av.
En tonåring och en yngre unge pratar vid en sammankomst i en park
En kvinna går förbi en västlig vapenaffär.
En man i blå kostym med megafon som går framför till folk klädda i blå dräkter
Två män, en i svart, en i grönt och denim, på ett dansgolv.
Två män i klänningskjorta och hålla mikrofoner sjunga tillsammans.
En grupp människor festar inne i en byggnad.
Person i en rutig skjorta som står i en folkmassa framför ett band.
En man i svart väst som spelar trummor.
En grupp människor sjunger i en fest
Fyra män spelar instrument och sjunger.
En skidåkare rycker på sig bakifrån goggles hos en expert bara tecken medan snötäckta berg fyller himlen i bakgrunden.
Folk dansar inne i ett rum där det händer en liten konsert.
Bandmedlemmar som leker med trumma majoren lyfter upp trummorna för att attackera en annan medlem.
En gitarrist med svart hatt som uppträder på knäna.
Två kvinnor dansar tillsammans framför ett band och en banderoll som säger "Live in Concert".
En man dansar framför ett band.
En grupp på sju män uppträder på en scen med mikrofoner och gitarrer när flera unga män och kvinnor dansar och tittar på.
En musiker i svart hatt spelar tangentbord.
En man drar en vagn hög med föremål.
En brud och brudgummen dansar i receptionen.
En kvinna i vit skjorta står vid ingången till en etnisk varuaffär.
Människor från en utländsk by samlar resurser.
Tre människor från Mellanöstern går igenom ett gäng glasflaskor.
Kvinnor i sari undersöker ett diagram.
En svart man i hatt sitter i en stol i sanden och håller i ett nät.
En man är skinande klädesskor.
En svart man utan skjorta kör en vagnslast full med varor.
Indiska kvinnor diskuterar sin uppgift på en grusväg.
Tre damer med halsdukar runt huvudet som gräver upp smuts.
En grupp kvinnor fyller i lite pappersarbete.
En mörkhyad man med turban ser upp tillsammans med andra klädda i sina infödda kläder längs en grusväg.
Fyra personer står utanför det vita huset.
En storögd kille i en blå jacka håller en öl och står bredvid en kille som håller hans näsa.
En man försöker sälja frukt på en livlig gata.
Fem attraktiva kvinnor som bär svarta mini-kjolar och röda toppar lutar sig mot en röd bil.
En kvinna avslöjar sin mage medan hon håller i en öl.
Du har två pojkar som spelar fotboll med varandra som båda är ute efter bollen.
En man i en formell outfit grillar eller kanske städar sin grill.
Revelers deltar i den kinesiska nyårsparaden med fyrverkerier.
En flicka står och en annan sitter vid ett träd
En man som går nerför en trottoar med två hundar på koppel.
En naken person som står på en sten.
En ung kvinna i rosa skjorta sitter på en veranda och väver med en vävstol.
En kvinna kollar sin väska på ett café.
Två killar delar hörlurar och lyssnar på musik på en tunnelbana.
En pojke som klättrar uppför ett berg.
En man marscherar framför två linjer av människor i uniform.
En man på landsbygden som använder jordbruksliknande utrustning i en träskmiljö.
En glasblåsare formar en flaska med en ugn i bakgrunden.
Fyra män klädda i vita spela saxofoner inför en publik.
Folk står på balkongen och däcket på en båt.
En ung man med mohawk börjar jaywalka tvärs över gatan.
En kvinna sitter på en matta omgiven av röda frukter.
En grupp människor står runt en man som sitter vid en symaskin utanför.
En kvinna och en ung flicka äter sida vid sida.
Två damer går på gatan; en av dem bär en stor last.
En kvinna i rött spelar gitarr och sjunger medan par dansar.
En järnvägsarbetare som arbetar på rälsen.
En man förbereder sig för att ställa in sitt skott under poolen i en poolhall.
En gammal kvinna med en vagn full av matvaror.
En man i grå jacka som står på sidan av en gata.
Två unga pojkar engagerar varandra under en flagbollsmatch.
En man med blont hår ser ut som en kvinna i en garnerad kostym danser på scenen.
En man i glasögon pratar med en kvinna medan han handlar apelsinjuice.
En man arbetar i en gruva eller en grotta av något slag.
Servitrisen lägger tårtan på ett bord vid en sammankomst.
En äldre man som läser en tidning sittandes åt sidan några hushållsvaror av plast och färgburkar.
Fansen hejar medan rullskridskorna går förbi.
Man i solbränd skjorta och blå jeans gör en rygg flip med bara fötter
Jag tror på tatueringsmannen.
En man som målar väggmålningar på trottoaren.
En asiatisk man som lagar kött över en öppen grill.
En vit man som håller i en pappersskylt med lite mat i brun skjorta.
Fem pojkar med tröjor och kepsar spelar football utomhus.
En man använder en mopp, medan två andra män tittar från bakgrunden.
En man hoppar på en bro av sten nära ett berg.
En kvinna med svart huvtröja står nära en gammal rostig lastbil.
Vi måste tänka på det här och det är ditt fel.
En man, som bär en officiell jacka och hatt, lutar sig mot ett sken medan han läser en tidning.
Sex personer vandrar i ett snöigt landskap.
En kvinna med svart hår och en röd rutig förkläde som lagar mat.
Tre arbetare i gröna västar som tar en paus.
Här är en grupp människor som väntar utanför på att bröllopet ska vara över och börja det verkliga firandet.
En liten vit hund står på ett ben för att fånga en boll.
Människor som promenerar i ett stadsområde i en stor stad där det finns eftergifter.
En man rakar sig i spegeln på ett fånigt sätt.
Två män rider nerför gatan på en cykel bredvid en grå byggnad.
En liten flicka kramar en artist i en Stitch-dräkt.
En man som har en blå jacka och fiskar i en flod och pratar med sin vän utan tröja.
En kvinna i en blommad klänning som bär grönt.
En man i vit skjorta som spelar en vit gitarr på en scen.
Cheerleaders uppträder på en fotbollsplan.
En man med tatuering på armen spelar dragspel.
Tre pojkar hälsar när de navigerar i vattnet.
Sju personer cyklar på en sandig bana.
En kvinna sitter framför en dator.
Några personer med gröna kläder bär en stor personal som ser ut som ett kors.
En kvinna i brun hatt kramar ett barn.
En äldre man som sover på en tågvagn med reflektion av andra passagerare bredvid honom i fönstret.
Två flickor städar och en flicka beter sig som en dåre.
En kvinna i en grön burqa och solglasögon går längs trottoaren mellan en väg och ett stängsel medan du trycker på något.
Militären hälsar på barn som viftar med amerikanska flaggor.
En tjej i vit topp sitter vid poolen.
En man som bär en officiell gul skjorta tittar på trafiken.
En vit hund med en tröja på och en svart och brun hund vidrör näsor.
En grupp unga elever poserar framför ett tecken.
Två män är ombord på en fartbåt som sitter lugnt i vattnet.
En liten flicka som står i ett badrum och borstar tänderna.
En man i en spetsig kostym går nerför gatan och märker inte den udda affischen till vänster.
Två män i svarta jackor som sitter på objekt som pratar.
En man i en jacka arbetar ovanpå en trappa.
En volleybollspelare hoppar för att slå bollen.
En man lyfter upp en kvinna i dans som deras pos för en bild som tas.
En man leker med en bebis på ett däck.
Två äldre män och en äldre kvinna sitter runt ett bord medan de pratar.
En flicka i rosa klänning kliver försiktigt över en pöl.
Tre kvinnor som bär affärskläder står framför ett fönster.
Ett barn ler medan de håller en flagga medan andra sitter i bakgrunden.
Två hundar brottas på marken i snön.
En liten pojke flinchar som en hjort kysser honom på kinden.
Fyra män gör en presentation medan ungefär åtta personer lyssnar.
Folk i kappor tittar på ett spel.
Två kvinnor, en med barn i barnvagn, pratar framför ett stoppet tunnelbanetåg.
En man och en kvinna på en motorcykel."
Någon hängde högt på en tråd nära en stor metallstruktur.
En samling människor som tittar på andra människor som spelar några instrument.
En grupp musiker som uppträder är omringade av det offentliga tittandet.
En man går en vit hund i koppel i en parkmiljö.
Polisen ser folk på en strandpromenad nära stranden.
Två kvinnor går genom gatorna och spelar tuba och cello.
En grupp på tre pojkar spelar fotboll medan en vuxen man tittar på.
En manlig leverantör väntar på att kunderna ska beställa öl.
En man som bär turban på huvudet ligger på knä och ber på en matta.
En person har ett hjul av en buss medan han mixtrar runt hjulet väl.
En arbetare är på toppen av en telefonstolpe och arbetar på ledningarna.
En kvinna på en Segway står med några män i en publik.
En liten kille i brun och grå tröja som trycker på en manuell gräsklippare på en inhägnad gård.
Man leder trafiken som en telefonarbetare utför sitt arbete.
En man i grön skjorta står framför en monter som säljer en produkt.
Musikerna spelar för publiken.
En grupp människor som spelar ett sortiment av instrument medan de går nerför gatan.
En man som står i vattnet.
En vuxen med ett spädbarn fastspänd på bröstpromenader i skogen med ett annat barn i bärgning
Ett marschband som spelar för publiken i en parad.
Marschbandsmedlemmar klädda i svart och blått spelar trummor och andra instrument.
En kvinna håller en svart skylt på ett gatumöte.
En ung dreadlockad kvinna står på scen, sjunger och spelar akustisk gitarr.
En grupp människor är i en skåpbil.
En grupp sjömän går längs en trottoar i en linje.
En ung pojke med baseballkläder som gör sig redo att kasta en boll.
En fågel flyger genom luften medan barnen leker på stranden.
En man kör en bår full av medicinska förnödenheter.
En man sitter i sin bil, med armen vilande på dörren.
Den bruna hunden har ett föremål i munnen.
En gatuförsäljare tenderar till sin monter med massor av barn leksaker och föremål.
En man och en kvinna sjunger på en scen.
En kvinna med mörkt hår och en blond kvinna i baddräkt har cocktails på en uteplats.
En ung pojke i skolan använder sax för att klippa papper.
En man som inte har en tröja och dansar ensam med slutna ögon.
En tjej i svart skjorta som spelar karnevalspel.
En man står i snön när solen går ner.
Ung muskulös afroamerikansk man, som städar en fisk, utan tröja.
Två svarta pojkar sitter i fiskebåtar med sina kastnät.
En ung blond pojke som borstar tänderna framför en spegel.
En man och kvinna i mellanösterländsk klänning springer nerför en gata.
En lycklig man i en blå krageskjorta skriver på sin dator.
Två svarta pudlar betslar lekfullt på en gräsbevuxen, manikyrerad gräsmatta.
En man som bär en läskig mask i en show.
Pojke går förbi mannen i orange overall som sopar sopor från gatan.
Vit man som sitter vid bordet med en dryck.
En ung man i röd skjorta gör tricks med en skateboard.
En liten pojke och en liten flicka på en veranda tittar på något.
En man i solbränd hatt sitter bredvid grön buskage och tittar ut över vatten.
En tonåring med randiga ärmar som spelar gitarr.
Fem unga kvinnor samlas i ett rum med gröna och blå stolar.
Två arbetare som jobbar på att sätta upp lyktor.
En man med mustasch och turban runt huvudet ligger i ett träd med ett verktyg.
Två mörkhyade män, en av dem med kniv, står framför något lövverk.
Medan solen går ner blåser pojken bubblor av klipporna nya sjön eller havet.
En man i grå strumpa tänder en cigarett medan han håller i en pop.
En man och en kvinna i orange trasa går längs en grusväg.
En schäfer hoppar i luften.
Fem personer står under en tältliknande struktur och firar den 25:e årliga Longboard Classic.
En kvinna blåser torka en ung pojkes hår i en hårsalong.
Asiatisk man i orange kostym och med glasögon som undersöker en ung flicka.
Äldre vit man som röker en cigarr
En man och en kvinna står vid en gatuförsäljares matstånd.
Två män står under ett vattenfall.
Dessa elever i klassen sitter ner och gör arbete.
En liten pojke med ryggsäck närmar sig en stenbåge.
Ett ungt par, både blond, kvinna i röd rutig jacka, bär en designer tote, bär bruna stövlar, korsar en upptagen stad gata.
Komisk man som trycker sin knytnäve mot en trasig betongpanna.
En man sitter på sidan av en trottoar med ett papper i händerna.
Asiatisk man i färgglada kläder skriva på sitt traditionella språk.
Två tjejer sitter i bruna stolar med drycker på bordet.
En man solar bredvid en pool med en vattenfallsfontän.
När man tittar ner från toppen av en klippa, klättrar en man upp på klippväggen i ett försök att ta sig upp till toppen.
Barnen är fokuserade på det grå objektet.
En man är klädd i vit peruk och skägg och lila klädnad och många människor tittar och tar bilder.
En äldre man och kvinnor som äter middag
Tre personer tittar på skulpturer gjorda av stenar belägna på en vattenförekomst.
Fotbollsspelare är uppradade på planen.
Slappna av under hyddan när någon går förbi med en fruktskålshatt.
En fotbollssparkare försöker göra ett field goal.
En fotbollsspelare tittar ner på en fotboll under en pjäs.
En fashionabel svart kvinna sitter på ett tåg.
En kvinna och en ung flicka går längs en vägg med siffrorna nittiosex prydda på den.
En grupp killar är inte han fotbollsplan spelar fotboll.
En kvinna med en röd ärmlös skjorta med svarta shorts springer.
En kvinna klädd i lager som tar hand om åkermark.
Två brandmän sprutar vatten från en svart slang.
En konstig pojke njuter av att röra vid höet.
Etnisk kvinna i traditionella kläder som sitter på marken genom konstverk i krita.
En person går på nattgatan under neonljus.
En man i ett vitt förkläde och handskar som stukar kol under en stor eldsvåda framför en trähög.
Sex personer verkar plantera något i marken.
En kvinna springer nerför gatan i ett maraton.
En gatuartist klädd som pirat offentligt.
Den här mannen åker skidor i den vita snön och går genom en kurs av något slag.
En affär på gatan som säljer grönsaker.
En rumpled man bär en bunt stockar framför en djungel.
En grupp afrikaner som flyr från något.
En asiatisk man och kvinna sitter ett bord, mannen på en laptop och kvinnan med en mugg.
En man som bär mask i ett rörigt rum.
Ett ungt köp som sparkar in sin karategi bredvid ett annat barn.
En man blickar uppåt medan andra tittar på honom på en stadsgata.
Rodeo repare på ett hus, försöker använda ett rosa rep, att fånga en ung tjur med horn.
Skådespelare poserar på ett evenemang.
Fiskare på marknaden väger sin fångst i slutet av en lång dag.
En kvinna med brunt hår som håller i en låda med ett snidat ansikte på.
Tre personer på en flygplats väntar på ett flyg
En man stryker tyget medan han röker en cigarett.
En indian i en senapsjacka skyfflar mycket snö.
En man i grön tröja har en rund, dekorativ kudde.
Folk på gatan kommer för att kolla kvinnobordet.
En flicka i randig blus sitter på en bänk nära en telefonautomat.
Två barn sitter medan en står över dem.
En pojke i gul jacka som håller i en röd gryta.
2 små flickor tecknar medan de lyssnar på ett band spela på en bar eller restaurang.
Två män pratar som fyra barn som springer förbi.
En kvinna och en man som pekar åt vänster står på ett gathörn framför en grön affär som säljer tobak och tidskrifter.
En man i en hård hatt tittar upp på något.
En äldre kvinna plockar upp en trädgren från sin stenveranda.
En arbetare som sysslar med vattenbesprutning överallt.
En orientalisk man med glasögon och en färgglad väst går nerför gatan med en tjej med blont hår.
En massa människor som pratar på en bar.
Yngre barn sitter och ligger på marken runt kläder och skräp.
En man i en rutig skjorta som spelar gitarr.
En leende flicka med en tatuering på handleden ligger ner i det vackra, gröna gräset.
En kvinna visar sina fingrar fulla av ringar i spegeln.
En kvinna i en vit och beige-strippad tröja svarar i telefon på ett kontor.
Två äldre män presenterar foton och diskuterar sina liv.
En man i röd skjorta och randig skjorta som sjunger var och en med mikrofon.
En far och son börjar en fisketur i en båt.
Två män i kostym sitter framför en publik medan en mans bild visas på en projektorskärm.
Folk pratar med en stor TV
En hund är på väg att få en boll som är på orange mattan.
Blond kvinna tittar ner över en träskena.
En man i arbetskläder och en vit hatt dränkt i vatten.
En kvinna visar känslor på en mikrofon.
En man med mössa lutar sig mot fönstret och läser en tidning.
Ett barn i gul skjorta klättrar upp i ett träd.
En tjej i gul t-shirt hoppar på ett fält en klar dag.
En man städar gatorna framför ett inhägnat hem.
Kvinnan i svart klänning håller ett papper i händerna när hon pratar in i en mikrofon.
En kvinna och två män spelar stränginstrument.
En man ligger på en fullsatt gata medan folk går förbi omedvetna om honom.
En man som hänger ut genom fönstret på ett tåg med svart jacka och hatt.
Tre barn rullar nerför en grön bergssluttning mot en parkeringsplats där en kvinna sätter sig i en vit bil.
Två skugglika figurer som står under en bro, två burkar vid deras fötter.
Kvinnor i färgglada utländska kläder talar på en marknad bredvid ett brödstånd.
Unga företagare som ger en presentation med hjälp av två bärbara Macbook.
En skjortlös man använder en rulle för att måla taket vitt.
Två unga flickor i skelettdräkter fastsatta i koppel.
En person i uniform står framför en tullbro.
Två äldre män sitter mot en blå vägg med sina käppar.
Folk sitter på stolar i ett rum med en person stående.
Två män klädda i vita skjortor står på en fest.
Ser ut som en man som transporterar en familj, bestående av en mor, en far och en son, till någon destination
En man sitter med huvudet nere på en tunnelbana.
Pojken i den svarta och gula masken pratar med mannen i den blå skjortan.
En kvinna stryker i sitt hem.
En man som sitter i ett tåg, tror att han är en dirigent.
Bilar parkerade på gatan på natten.
En militär man går framför en procession av människor under en parad.
En kvinna som försöker skapa en isskrift.
Två män med svarta skjortor sitter bakom sina egna färgglada trumset.
Tre flickor står utanför, en flicka gråter.
Bandet uppträder på fotbollsplanen.
En grupp byggnadsarbetare går.
Simmare gör varv i en pool.
Två fotbollslag tävlar i en fotbollsmatch utanför.
En manlig och kvinnlig kock vakar över köttet och majsen de lagar.
Två barn äter glass på en bänk.
En man med skägg sitter med en gitarr som har öppnat sig, och trådar exponeras.
Ett par sitter tillsammans och tittar på en bildskärm.
En man spelar en speciell gitarr och tittar på en TV.
En byggnadsarbetare vilar en stund.
En man med gitarr har trådar på fingrarna för att spåra deras rörelse.
En kvinna som tittar på en mans datorskärm.
Två personer kommunicerar medan de sitter på en bar.
Några poliser på en scen.
Två poliser på ett förortshem som filmar ett polisområde med gul tejp.
Två personer i kostym går upp.
Ett barn står på en gångväg med solen mot ryggen.
En man som spelar gitarr och en kvinna som bär handske.
Två muslimska män sitter på sitt bås för att tjäna lite pengar med den verksamheten.
En svart man som bär en stickad hatt mönstrad med snöflingor ler något.
En äldre man som sitter på en fällstol och tittar ut på gatan.
Man arbetar på beige snideri medan bär gula öronskydd.
Den vita och bruna hunden hoppar upp i luften, ovanför snötäckt mark.
Folk som står runt en svagt upplyst bar och umgås.
En liten grupp tonåringar går längs en gata tillsammans klädda med handgester och med strumpbyxor och minikjolar.
En asiatisk dam i en röd jacka som tar ett foto
Folk i kostym värmer upp framför en brand.
Ett par poserar för en bild på fältet.
Tre pojkar kämpar med varandra och sträcker sig efter en påse skräp.
Ett äldre par som ler medan de står framför en stor byggnad.
En man som bär huvudduk och ländduk lägger och jämnar ut en asfaltyta nära en skog en varm dag.
En gentleman som använder en fackla för att försegla en löpare till en galla.
En man använder en blåslampa på ett provrör medan eleverna tittar på i bakgrunden.
Ett barn som visar det är mycket trött och sömnig.
En hiss i ett köpcentrum ligger framför en gul och grön vägg.
En person klädd i rött och svart utanför en sprucken vägg.
Ett barn står vid en pool med en stolpe för att rensa poolen.
En pojke med en blå t-shirt som ligger på en säng.
En man med glasögon tar en bild av ett tåg.
Tre tonåringar pratar nära en vägg.
Många människor i ett rum fyllt med halloween dekorationer.
Kvinnan på mobilen springer i snön.
En svart man som pratar med en kvinna på gatan.
Två personer tittar ut genom fönstret och tittar på radarn.
Personen i den blå skjortan och den blå hatten rider på en vit häst.
En far lagar frukost med sin dotter.
En ung pojke är ögonbindel med en mask och slår en pinata medan en ung kvinna och småbarn klocka.
Två män pratar medan de sitter på en parkbänk.
Två pojkar springer runt en tjej som ligger under ett paraply.
En byggkille med sin hatt på pratar i telefon.
En person kör över en torr terräng på ett All Terrain Vehicle, bär mestadels grön växel.
En man som har spikar på ett skjul.
En man klättrar upp på sidan av ett berg.
Två personer klättrar.
En blond klättrare med en vit skjorta skalar en stenklippa.
En man i en limegrön väst styr trafiken
Två personer i regnutrustning är löv som blåser i gräset under en regndag.
En man som bär glasögon rakar sig i en spegel.
Många män i gula skjortor och en kvinna i orange skjorta tar en spinklass och ler.
En man i grön skjorta går en spinningskurs.
Två damer ena med fingrarna i fickan och den andra med en drink i handen på en fest.
Damen gör en gymnastisk rörelse medan böjer sig bakåt och håller ett lila band.
En banddansare hoppar genom luften med huvudet tillbaka under en tävling, grönt band bakom henne.
En maskerad kvinna med glasögon håller i ett barn.
En hona i gult bär en kirurgisk mask håller ett spädbarn.
En gul ballong flyter över en stenbyggnad.
En liten flicka i röd rock med en korg på sidan.
Kvinnor som pratar medan de väntar på något.
En kvinna serverar mat vid vägkanten.
En man med gul väst fungerar på gatan.
En liten grupp människor, däribland en cyklist, förbereder sig för att korsa en gata i staden.
En leende vandrare poserar på toppen av ett snötäckt berg
En man på en ATV med två barn på baksidan.
Pojke sitter och tittar genom ett glasfönster på en tågstation.
En person i en utstuderad mask håller upp en fackla framför en folkmassa.
Två personer spelar ett spel i en arkad.
En man i rullstol knuffar längs stranden medan två barn leker i förgrunden.
En jockey klättrar en ramp bakom sin häst.
En man, i en gul keps och solglasögon, är ombord på någon sorts båt på vattnet.
Fyra män flyter i en blå båt medan boskap betar i närheten.
En liten flicka i grön rock och en pojke som håller i en röd släde går i snön.
Infödda amerikaner utför en traditionell dans eller ceremoni.
Två personer står framför en tegeltågsstation och väntar på ett tåg.
Pojke står nära tvätten hängandes för att torka.
En pojke försöker sig på skateboarden i parken.
En man i en grön huvtröja försöker göra ett trick på sin skateboard i en park.
Fem unga kaukasiska vuxna tillagar mat tillsammans i en matsal.
En ukrainsk man i kostym utför en dans på scenen.
Ett par i traditionell holländsk klänning dansar på en festival.
En festival pågår på gatorna.
En man som kliar sig i armen medan en flicka sitter vid ett bord.
Tre män samlas runt ett fruktstånd.
Två killar på stranden som leker i sanden, med en vän som försöker sparka den andra.
Ett par och deras barn slappnar av på en kamrat.
En man i röd skjorta som klättrar på en klippa med sina bara händer.
Arbetare på Starbucks restaurang visar upp sina lokaler.
En man i vit t-shirt och jeans använder en skiftnyckel.
Tre personer i kostym går på trottoaren.
En man som bär en knapp-up skjorta spelar en flöjt medan han bär en flaska och en stor pinne med många flöjter i ena änden.
Två pojkar i blå tröjor omfamnar en bild.
Sex personer på scenen gör sig redo att buga.
En hund med munnen öppen för att fånga den röda bollen.
Äldre kvinna som sitter i en kaninbur med två vita kaniner i knät.
En brud och brudgum som skär sin tårta.
En kvinna går mot en vaktmästare som bär regnrock och trycker på en städvagn.
2 svarta flickor i lila skjortor sitter nära ett grönt staket.
Svarta skolpojkar i uniformer gör affärer med en vit man under garagedörren.
Vissa väntar i kön.
En tjej i kattdräkt tittar på en bok.
En kille i gul och lila dräkt som hoppar från en trappa.
En gammal kvinna klädd för kallt väder i hatt och solbränna rock med en käpp som håller en liten bit papper.
Folk springer i ett lopp på en gata.
Runners i olika färger kör vänster på foto, med man i framkant viftar på kameran.
Gammal kvinna på vintern går förbi en glamourbutik.
En tjej i en ljus utstyrsel leker i löven.
En grupp löpare avbildas när de springer ett maratonlopp.
En del människor vilar nära en skog och nära en flod.
Från en tjej som tar itu med en annan, säger jag håll fast vid din drink!
En judisk man håller huvudet av en annan man som har böjt sig ner mot honom.
En man och kvinnor som går förbi ett varningstecken.
Två små barn ligger på en veranda i sovsäckar.
Människor i klungor av tvåor och treor står runt en fontän utomhus.
Två äldre män samtalar stående i en gammaldags, asfalterad gränd som gränsar till färgglada byggnader.
En person som bär en gul skjorta går nerför gatan och bär en stor korg.
En man och en kvinna sitter på en bänk och läser böcker.
Runners tävlar förbi medan en skara åskådare tittar.
En stor grupp människor kör ett maraton och övervakas av åskådare.
En grupp simmare dyker ner i en simbassäng.
Framslags simning ras repade bort varv områden.
En idrottsman som simmar under ett simmöte.
En man i svart skjorta som håller upp ett papper fullt av matematiska ekvationer.
Fem vandrare går nerför bergssluttningen.
En man är ute på en sko skinande stå skinande en kunder skor.
En man med hörlurar blandar musik.
En man i vit skjorta lutar sig över en dator.
Fem män i ett laboratorium tittar genom mikroskop.
En vietnamesisk man som kör en traktor genom en ravin medan en kvinna rider på baksidan.
En kvinna med en blå skjorta som skriver på en laptop.
En trumma hammar rasande ut anteckningar på sina instrument när han spelar på scenen.
En man med en svart skjorta som sjunger in i en mikrofon.
En man leker med sin skateboard på en gata.
Två ungdomar tittar på en fontän.
Två män använder skateboard mitt på gatan.
En man skateboardar medan två andra tittar på.
Två manliga bandmedlemmar spelar gitarr framför en mikrofon.
En man som lagar mat i ett kök.
En gammal man och två barn är på verandan och tittar över räcket
En blomsterförsäljare på trottoaren som förbereder sig för att skanna en kunds köp.
Ett barn ler mot en kvinna på andra sidan bordet.
En präst sitter i en gammaldags träbekännelse.
En hund i vatten med huvudet tuppat åt sidan tittar på en boll.
Två ljust klädda kvinnor med hattar tittar på något.
En man med kort hår och skägg håller ett barn.
En ung man som tittar på rått kött hängande.
Cyklist går cykel nerför en tunnel som inte tillåter cykling.
En flicka med skyddsglasögon ler mot kameran.
En medelålders man bär karatedräkt medan han övar med en annan maskerad individ.
Mannen och hans slädhundar färdas längs en snöig väg.
En ung pojke i blått leker i ett rum med många leksaker.
Slumpmässiga människor på en flygplats som gör olika saker.
Den svarta och bruna hunden springer med något i munnen.
En vit hund med flytväst följer med en man i en båt.
En stor grupp kvinnor, som bär rosa skjortor och svarta byxor, har armarna upplyfta med höger arm utsträckt och vänster arm böjd inåt.
En man tittar på en kvinna när hon cyklar förbi honom.
Två män tittar på framsidan av en snöskopa maskin.
Ett barn som bär kappa ser tillbaka på någon.
En grupp kvinnor står nära en grupp armémän.
En man och en kvinna för en diskussion medan militära medlemmar ser på.
En grupp barn som står i en cirkel och håller varandras händer.
Soldater i uniform stirrar på två små barn.
Två män i militäruniform står framför en lastbil med leksaker.
En kvinna som håller ett litet barn med tummen upp.
Soldaten tittar på digitalkameran som ett barn med juice box tittar på honom genom nyanser.
Två män i militären och en pojke poserar för en bild.
Soldater står i formation utanför en byggnad, och en man klädd i gatukläder står nära dem.
En grupp bybor förbereder sig för en regnstorm.
En man i militär kamouflage och en mörkgrön hård hatt håller ett inramat barns krita teckning.
En arbetare i en hård hatt blir intervjuad.
Män knäböjer runt ett brädspel utanför på en kaklad yta.
På den här bilden ser vi en man som lagar mat i ett kök.
En äldre kvinna sitter i bur med två bruna och vita kaniner.
En man skyfflar snö mellan två svarta fordon.
En hane som åker skateboard nerför en trottoar med en vit randig skjorta och svarta byxor.
En äldre man som cyklade med en stor vit byggnad bakom sig.
Bald man i en skjorta en slips som står runt mat och dricka vin.
En fotbollsmatch spelas av lag i blått och rött.
Den här mannen bär en röd hjälm och flip-flops och kör en Spyder.
En kapten kollar sina passagerares livvästar.
Två kvinnor ler och pratar med varandra medan de båda håller en burk öl.
En man med upplyft hand.
En grupp människor samlas för en måltid i business casual klädsel.
En man på en smutscykel i luften tävlar.
En utomhus cykel händelse med Braun markeringar på väggarna, en cyklist kör har gått fel med sin cykel flyger upp i luften medan andra tittar.
Här är en gråtande bebis som hålls fången av sin mormor.
En man i mörk tröja sitter vid ett bord med en röd penna och en tidning.
En flicka som rider en ponny med flätor och rosa rosetter
En man med skägg och svart skjorta som tittar på ett kuvert på ett kontor.
En kille använder en bulldozer, och de arbetar på avloppsledningarna.
En grävsko gräver en dike utanför en byggnad.
En kille som står vid en elstolpe och poserar på jobbet.
En man som bär brun rock och latexhandskar tittar på något i fjärran.
En hane med hatt och glasögon står runt omkring.
Ett par i svarta rockar tittar på kameran med trevliga uttryck på sina ansikten.
Ett par är förblindade av ljuset från en kamera.
Två personer sitter på en bänk med utsikt över en stor mängd fönster.
Vid en militär ceremoni deltar pojkscouter.
En man i en tröja poserar i sin vikinghjälm medan en annan man i en rock tar en bild med sin kamera.
En man i rutig jacka arbetar med blommor.
En man och en kvinna håller hand på ett gräsfält.
En man sitter på trottoaren bredvid sin skoputsningsstation.
En grupp scouter står i en alert position.
Krigsveteraner deltar i en minnesceremoni utomhus.
Ett gammalt par med sina vinterjackor står framför ett köpcentrum.
Utländska militanter eller myndigheter som upprätthåller fred och ordning på en gata i grannskapet.
Kvinnan cupping vatten med händerna över badrum handfat som barn står bredvid henne.
Två män står framför en solbränd byggnad.
En person observerar två personer som sitter på en tegelbänk och tittar igenom föremål som tagits från en gul hink.
En man med vitt hår som går längs trottoaren.
En grupp unga etniska barn som utför en dans i traditionella färgglada kläder.
Kvinna stretching i ett kök medan blanda ingredienser i en skål.
Två vuxna är ute och pratar, medan en liten pojke tittar på dem.
En man försöker titta på sin TV på en offentlig plats
En man som sover medan han sitter på en buss med väskan i knät.
Gamle man som spelar saxofon på gatan.
En kvinna sitter i en brun stol mitt i ett köpcentrum.
En kvinna som målar en annan kvinnas naglar är ljuslila.
En ceremoni med en man som talar och en annan man som justerar dräkterna på en annan person vars ansikten delvis är täckta och hålls i en moské med många iakttagare.
En mogen asiatisk man står i en grå hall.
Två fotbollsspelare, en i vitt, den andra i maroon, spelar och spelaren i vitt är ute efter en rubrik.
Man går förbi en busshållplats med graffiti.
En man i blå skjorta med mustasch som pratar på en mobiltelefon
Den ena konstruktören lägger sig för att vila medan den andra sitter i en stol.
I bakgrunden finns det 3 personer på stranden bland flera kanoter, och den unge mannen i förgrunden paddlar genom vattnet, samtidigt som han bär flytväst och ler.
Lägerledare samlar och organiserar information och unga flickor för sin lägergrupp.
Två män, den ene yngre och den andre äldre, var stationerade på vad som ser ut som en kontrollpanel på en flygplats.
En skara människor deltar i ett utomhusevenemang.
En kvinna klädd i rosa håller en bok framför ett veteranminne.
En liten flicka sticker ut handen för att ge maratonlöpare en high-five
En grupp barn och vuxna som alla bär blå ryggsäckar står på en trottoarstig i öknen.
En man knäböjer på en brygga medan en hund hoppar i vattnet bredvid honom.
En hund med en glänsande hund taggar ändrar kurs på hans steg
En massa människor på restaurang äter.
En liten pojke i en grön och vit uniform springer mot en röd, svart och guldfotboll.
En man står utanför glasdörrarna på ett konstcentrum.
Ett litet barn med munnen vidöppen för en stor sked mat.
Svart kvinna i orange klänning skyfflar korn.
Kvinnor i Saris går längs en grusväg.
En man sitter vid ett stökigt datorbord i ett vitt rum.
Två män står på vägen, det verkar nästan vara någon sorts film som spelas in en solig dag i Kalifornien.
En grupp människor står utanför en byggnad.
Ungt barn slappnar av och njuter av ett mellanmål medan hon sitter i ett badkar med fötterna ut.
Människor på en marknad som köper frukt och grönsaker
Det är en livlig gata i Indien där det finns affärer och människor går, cyklar och gör sina dagliga ärenden.
Den lille pojken har sett fotografen från ovan.
En kvinna och hennes barn rullar ett mindre barn i en barnvagn på en tegelstig.
En liten pojke med blå shorts och gul skjorta trycker på en barnvagn.
En man i röd tröja pratar med en grupp barn i skogen.
En blond artist står på scen i en vit outfit.
En man håller i en fiol medan han sjunger in i en mikrofon.
Två blonda damer sitter på en soffa och dricker vin.
En man med blå jeans och väst ligger på en stadsbänk bredvid en ölflaska.
Flera små barn spelar basket.
En ung vit man som bär glasögon rakar skägget med en elektrisk rakhyvel.
En kock som kryddar nybakade popcorn vid fönstret.
En man i röd jacka med snöutrustning är mitt uppe på en snowboard med en röd struktur i bakgrunden.
En sångare uppträder på scen på en konsert.
En man med tatueringar står mitt i en scen klädd i vita byxor medan tre andra står framför honom.
En ung kvinna balanserar på en upphöjd plattform.
En man i mörka badbyxor leker med en pojke i röda badbyxor på stranden.
En afrikansk man som sitter på en bänk ritar en bild.
En kvinna i svart rock sminkar sig i ett tåg.
En kock som lagar lunch i köket.
Två pojkar tänker på vad de vill köpa och två pojkar hämtar pengar de tappat.
Tre kvinnor i jackor korsar gatan.
En kille hoppar i luften medan en grupp människor står och ignorerar honom.
Den lilla bruna hunden hoppar över tegelväggen.
Någon går längs en ensam väg i en nästan övergiven gång.
En kille som mediterar på gräs med slutna ögon
En man i en keps skapar en skulptur av en man.
Två män med vita skjortor och slipsar dricker.
En man i en grön och vit randig skjorta bär en stor korg på axeln.
En kvinna som bär rött talar genom en megafon medan hon går framför en banderoll.
Unga flickor väver majsstjälkar till genomtänkta mönster.
Folk äter mat i en livlig restaurang.
En kvinna korsar gatan, kamerans utsikt är mellan två bussar.
En publik tittar på två sittande musiker och en talare som står på ett podi.
Två dansare, en man, en kvinna, gör en rutin i en dansstudio.
Många kvinnor dansar på ett brunt dansgolv
En brun bil dyker nerför gatan, medan folk går över hörnet.
Folk är trånga runt en förfallen buss på gatan hörnet
En man i blå shorts och en man i telle och orange shorts skördar en bale.
En man i tröja viftar med flaggor.
En man i gul kostym klättrar över ett trasigt staket medan en annan man tittar på.
En kvinna går framför en filmreklam.
Några ungar samlar löv och lägger dem i sopsäckar.
En man som ger en presentation framför en projicerad bild.
En man, som bär en kostym med en namnbricka, talar i en mikrofon, medan han står framför en videopresentation.
Cowboy rider en häst i en parad som åskådare klocka från trottoarkanten.
Tre unga män samlades vid ett bord och drack och diskuterade.
Två kvinnor med paraplyer springer tvärs över gatan i regnet.
En fastare som bär hatt blir fotograferad.
Ett par skär tårtan med en publik.
En kvinna och en hund är i ett fält av starkt grönt gräs och lysande blå himmel.
En mellanösterländsk kille som säljer saker på gatan.
Tre män i matchande reflekterande uniformer samlas framför en dekorerad vägg.
Folk på trottoaren försöker skydda sig mot regnet med paraplyer och en tidning.
En kille och flicka på klippor som fiskar i en vattensamling.
Mannen i en nålstickad jacka arbetar med ett föremål.
En liten pojke prestends att slå en annan unge i templet medan de äter lunch.
En man som målar en golvblå med bara byxor och hatt.
En pojke håller en blå pinne, medan en man håller en pinata ovanför honom.
Två hundar leker med en boll i snön.
Ett barn undersöker en bit sten genom ett förstoringsglas.
En man i grå skjorta har sina armar upplyfta.
En pojke surfar på en gul tavla över den ljusa blå vågen.
En man som grimaserar medan han använder en motoriserad tandborste.
Två pojkar, en klädd i en röd Chiefs tröja, leker nära en strand.
Två små barn leker.
En indian med saknade tänder, en röd hatt och en röd vinge eller filt ler.
Flera kunder handlar grönsaker på en bondes marknad.
En California Golden Bear quarterback faller till marken efter att han kastar bollen till sin mottagare som jagas av Stanford försvar.
Människan går sin hund över intressant yta.
En liten flicka äter en korv med handen.
Två män i svart springer genom en skog.
En stor folkmassa som sitter vid bord i ett stort tält.
Ett barn tittar uppmärksamt när en kvinna använder en MacBook laptop.
En man tar en promenad med sin hund under solnedgången.
Män som bär färgglada jackor finns runt en landad helikopter.
Två äldre kvinnor sitter i stolar och pratar med varandra.
Fyra människor skördar på ett fält.
En man och en kvinna står tillsammans när hon röker en cigarett.
En servitris på en restaurang städar ett bord.
En man i blå jersey och blå keps tillagar mat medan han står vid en disk framför ett fönster.
En man med ryggsäck går nerför en pir bredvid vattnet
En ung kvinna med svart hår och långa vita stövlar poserar i en kort klänning med vit bakgrund.
En pojke med gitarr sover bredvid en betongstruktur.
Asiatisk kvinna spelar musik inne i en tunnelbanestation.
En grupp människor pratar och äter.
En man spelar en orgelkvarn med en leksaksfågel i en bur.
Brandmän släcker en brand i en husvagn.
En person i svart skjorta lastar av föremål från en lastbil.
En kvinna i svartvit klänning som leder en kör.
En man som spelar flöjt framför en blond kvinna
Ett lokalt band har en spelning i en hall
En man står med slutna ögon och röker en cigarett.
En man utan tröja hoppar av en avsats i vattnet.
En skäggig man som bär en bast arbetar med ett projekt med eld.
En skjortlös pojke i flip-flops kör en wheelie på sin cykel.
Män i röda byxor marscherar med pinnar i sina händer och starkt ljus går runt dem.
En del människor väntar på en trottoar för färsk mat.
En ung flicka i lila jeans och en lila jacka står på armar och ben med ryggen mot marken.
En man i svart hatt med grön rand spelar dragspel.
En kvinna i solskyddsrock sover på en man med glasögon.
Hockeyspelare och domare förbereder sig för en face-off.
Män sitter vid ett bord med namnskyltar och framför en stor skylt.
En stor grupp människor tittar uppåt.
Fyra skäggiga män sitter i en restaurang och ler mot kameran.
Flera jakthundar samlades som en publik klockor.
Två kvinnor i ljusblå skjortor lägger en stenpanna i en trädgård.
En man som liftar med en påse har kommit tillbaka.
En grupp människor går på en stig genom skogen.
En skäggig man ger gester med händerna i köket.
En man i ett blåkontrollerat förkläde använder rengöringsmedel för att sanera en yta.
En vaktmästare moppar trägolvet i ett klassrum.
En man med långt hår spelar gitarr.
Två hockeyspelare väntar på att en puck ska släppas av en domare.
En person i vit t-shirt hoppar framför en sjö.
Barnet använder ätpinnar på välte köksföremål.
Unge man klipper sig av en annan ung man.
Svart man bär Run DMC t-shirt ger en annan svart man en frisyr
Tre män samlas runt medan en styr en kamera.
Den svarta pojken i den grå t-shirten skakar sina händer.
Man utanför i regnet främjar en 50 % rabatt försäljning.
Unga kvinnor i färgglada dräkter höjer händerna i lycka.
En man i grå skjorta får håret gjort med folk som står runt honom.
Ett upplopp bryter ut på gatorna i en asiatisk stad.
En tjej i randiga strumpor sover på en grön soffa med röda kuddar.
En soldat och hans dotter bjuder på lunch.
En man i grå skjorta klipper sig.
En pojke får sin frisyr av en annan pojke med vänner som tittar.
En man i vit skjorta klipper en annan mans hår.
En man står nära en pool med sin grå skjorta delvis över huvudet.
En ung flicka i rosa leker med en rosa leksak på asfalt.
En man står på ett metalltak och sprutar röd vattenslang.
En hund står i snön och tittar på kameran
En man sover ute på sten.
Det är många som handlar i klädaffären som säljer Carhartt.
En flicka i rött och en man i svart dans
En skäggig man med dreadlocks i en orange skjorta har stamansiktsfärg.
En man som läser en sen nattbok på soffan.
En liten flicka som hoppar upp för att landa på en gul cirkel vid en stänkplatta.
Ett barn som dyker in i en allmän inomhuspool.
En kvinna i svart och solbränd jacka, solbränd hatt och röda byxor har precis satt en golfboll.
En person som fotograferar utanför i snön.
En man i en hiss tittar på spegeln på väggen.
Kvinnan bär en strumpa, står i en tunnelbanetunnel.
En svart gitarrist i en gul träningsoverall och svart fedora sitter på en offentlig bänk och spelar gitarr.
Tre damer med tyg som tittar på en telefon.
Smickrande småbarn som bär en blå skjorta ler medan de sitter på en gungställning.
Flickor i knäskydd och rullskridskor står tillsammans.
En grupp människor i vildmarken som packar lådor fulla med mat.
Kinesiska medborgare går genom torget.
Fotgängare promenerar omkring i ett torg framför en stor byggnad.
En kvinna i blå skjorta sitter på trottoarkanten.
En man som vänder sig om och ler när han går nerför en livlig gata på natten.
En dam som bär på mat över en bro.
Pilot i cockpit i en grön väst på väg att slå på en strömbrytare.
En gammal man säljer frukt.
Två arbetare i hårda hattar arbetar på maskinen i närområdet med taggtråd.
En skäggig man visar upp vad han just lagade.
Män jobbar utomhus och man klättrar på något.
En ung pojke springer förbi en graffititäckt vägg.
En man med en stor växt läser en tidning om hur någon (förutom honom) är en idiot.
En familj i en timmerstuga ställer upp för en födelsedagsfest
En pojke som försöker övertala en flicka att följa med honom in i affären.
En man sjunger medan en rödhårig kvinna väntar på sin tur.
En man och kvinna i svart lämnar och går in i ett kök, kanske för en St Patricks dag fest.
Flera personer köper empanadas från en liten empanadasbutik.
Lumberjack i sin säkerhetsröda overall, blir snygg med sin orange hårda hatt när han skär ner träden.
Barn leker i en rondell.
En kvinna i gul skjorta dansar barfota på en blank yta framför skogsbruket.
Brandkåren är på plats för att hjälpa till vid en olycka.
Två män drar på ett nät nära stranden med vågor kraschar bakgrunden
Den här mannen sover på en bänk.
En man, som bär glasögon, är bergsklättring.
En gammal man och en gammal kvinna blåser upp en varmluftsballong.
En man i gul utstyrsel som ser några män spela schack.
En svarthårig man klipper sig.
En man står bakom en bar som serverar flera sorters öl.
En man sjunger med en clown bakom.
En kör klädd i svart uppträder för en publik.
Ett par gör sig redo att ta bröllopsfoton.
Fem personer i ett lopp går bredvid varandra.
Killen i vit fuzzy jacka spelar gitarr medan en man i lila knapp upp sjunger.
Fyra män på en fotbollsplan medan sprinklern är på.
En liten vit hund springer över ett gräsfält.
En man i uniform styr trafiken när folk korsar gatan i en korsning.
En vit vägg med bilder med en liten pojke som tittar på dem.
Två barn leker på vägen medan deras föräldrar väntar och sitter på bänken.
En fotbollsmatch ska börja.
Två kvinnor som går klädda i blått på ett fält.
En man i skotsk dräkt i en parad
Folk på någon typ av utomhusmässa.
Två pojkar pratar medan en sitter på en mula.
En städare i ett stycke moppar golvet framför sin trehjuling full av förnödenheter.
En skäggig man som njuter av ett varmt bad.
En liten flicka står på en kullerstensgata och tittar på bubblor.
Två personer i vita toppar och svarta förkläden.
En unge som försöker klättra upp och springa genom en skateboardbacke.
En liten flicka i jeans och en blå skjorta sitter på en gunga.
En kvinna som bär blå kläder visar en bildbok för flera små barn.
Barn sitter i stolar med musikstånd i bakgrunden.
En grupp barn som har fjärilsutskärningar i luften.
En kvinna i ett förkläde letar efter bröd.
Tre personer som bär livsvästar paddlar längs med en kanot på en liten flod i ett kärr.
En man klädd som 80-talsfilmen Batman.
En liten flicka i rosa står bredvid en liten blondin och tittar på kort.
Barnen står under ett paraply i en flod.
En grupp människor ser en man stå på en pall klädd i en stringtros.
En bedårande ung pojke roar sig.
En ung flicka i blått i en sväng utanför med slutna ögon och händerna av svingens kedjor.
En grupp människor står framför en matbil.
En grupp människor som sitter ner till en måltid i en gammal träbyggnad.
En man använder en kvast utanför en affär.
Pensionären, som bär träningsoverallen, åker skateboard genom parken.
Denna marknadsplats har flera leverantörer som säljer frukt, grönsaker och andra produkter.
Två barn njuter av bakverk medan de sitter i stolar bredvid varandra.
Personen som bär den röda hatten är på berget.
En man i svart skjorta tar av sig arbetshandskarna vid en röd grind vid en byggarbetsplats.
En ballongförsäljare står på gatan medan motorcyklar kör förbi.
En man i en bergig region arbetar med en cirkulär bit aluminium.
Två dykare fotograferar under vattnet tillsammans.
En ung pojke står bredvid ett öppet skåp, och han är täckt av mjöl.
Två små barn leker på en staty.
En kvinna som bär röd rock och randiga byxor lutar sig mot en man som bär svart hatt och röker en cigarett.
Två musiker i svart spelar saxofon och trumpet runt tallar.
Ett barn i rosa rock står mitt i en hög med tomma plastflaskor.
Här är en man som protesterar mot vatten på flaska.
Folk som går över vid ett stoppljus framför en stor byggnad.
En äldre kvinna kollar sin klocka.
Två kvinnor med hattar går ifrån varandra med sitt bagage.
En rullskridskor utför en tågrip från en böjd vägg.
Sex personer i vita hattar går på en gångväg täckt av snö.
Två personer joggar på en stig.
En person som bär ett vitt klädesplagg med en brun väst står bredvid en matta där en man ligger lutad bredvid vissa föremål.
En hund springer genom skogen.
En stolt far med sitt barn och sin hund sitter i en solstol utanför och tittar på sin son.
En man och en åsna som bär på halm går längs en väg.
Två knubbiga, medelålders kvinnor står på en parkeringsplats bredvid en tom kundvagn.
En kille hjälper en yngre tjej att klättra med träd i bakgrunden.
En rosa tjej dras upp med klättringsredskap av en man.
En vuxen manlig och kvinnlig balans på en såg.
En man sitter framför sin grå laptop.
En man och tre barn som cyklar med fyra säten.
En kvinna äter middag med sin hund när hon sitter på soffan och det finns fyra tända ljus på bordet.
Två små flickor tittar ut på flygfältet med förundran.
En man klädd som jultomten lämnar sin Prius framför Ruby's Diner.
Två unga flickor som leker ute på lekplatsen.
Folk åker skridskor på en upplyst plats nära en plats som säljer alkohol.
Fyra personer sitter vid ett bord och äter.
En ung pojke som bär en grå tröja målar på ett papper med kritor.
Mannen är en rosa skjorta som står på trottoaren.
En kvinna som sitter i baksätet på en SUV och lagar mat.
En person som sprider lim på sulan på en sko
Unga män och kvinnor som skriker med allvarliga ansiktsuttryck.
En man och en kvinna handlar i en stor järnaffär.
En man på en hög stege målar utsidan av ett hus.
En man som gör en midair kick på en karateturnering.
Två arbetare står på ett tak medan de reparerar en skorsten.
En kvinna som håller hand med ett barn som går på en bänk.
Ett nytt barn på sjukhuset, insvept i filt, sovande.
Två barn sitter på en stadion.
En brun och svart hund som springer på en strand nära stranden.
En skäggig man i grön rock stirrar in i kamerans lins.
En kvinna plockar majs, hälften gömd av stjälkarna.
Ett barn leker med sin fars stövlar.
Män kör bort från en brygga i en orange båt med en utombordsmotor.
Fyra män och en kvinna sjunger en sång på ett evenemang.
En far och hans barn väljer ut en julgran.
En grupp människor cyklar.
En liten pojke som sitter utanför och tittar på upplysta lyktor.
En tjej som sitter på en bänk.
Grupper av människor sitter på trappan med utsikt över trädgårdar och fontäner.
En av bandmedlemmarna som spelar hans trombon.
En hund springer vid stranden av en sjö, kulle i bakgrunden.
En lycklig pojke hoppar i sanden.
Två pojkar och en flicka som gör skolarbete i ett klassrum med en grön vägg i bakgrunden.
Ett barn sitter bakom ett konstgjort bord.
Waist ner bild av en surfare rider en liten våg.
En man som sitter på en grön stol på en flygplats.
En grupp människor i blandade åldrar sitter på en buss som har röda nackstöd.
En pojke och flicka står nära en clown.
En grupp människor sitter vid ett rundat bord inomhus och äter mat.
En hundvalp hoppar på en säng.
Ett barn sover på golvet med ett uppstoppat djur.
Gruppen väntar på resan.
Tre små flickor sitter vid ett rött bord med ett tomt grönt bord i bakgrunden.
En man som utför ett skateboardtrick, med gatlyktor och trafikljus bakom sig.
Män med svarta västar står där bak när en kvinna lyfter en gul flagga.
Två män av latinamerikansk härkomst arbetar vid träbrädorna.
Mannen i orange skjorta och skor står bland lådorna medan han håller en låda i handen.
En grupp män får sina bilder tagna i steg.
Två unga flickor i röda baddräkter som simmar i vattnet.
Flera hundar slåss i en gränd nära en silverbil.
Två män, en som håller i en mikrofon, talar medan de står på ett trägolv avsett för ett idrottsevenemang.
Två asiatiska kvinnor som surfar i en affär.
En pojke i röd skjorta klättrade upp på toppen av ett djungelgym medan andra barn leker längst ner.
Fyra personer tittar på en man som står i floden
En man står framför en tegelvägg med staden i bakgrunden.
En man klädd i juldräkt, med skägg och glasögon.
En ung kvinna med grå skjorta tittar på en brun keramikbit.
Man på toppen cykelstolpe sitter på cykel med en kall drink.
En man i vit skjorta ger detaljer till små skulpturer.
Olika människor ute och omkring på en offentlig plats på en höstdag.
En man täckt med en röd skjorta och solglasögon är avkopplande på en veranda med en tidning.
En man med tennisboll som leker med sin hund.
En professor håller en föreläsning för elever i ett klassrum.
En kvinna gör en lerkruka.
En man med hatt och blå jacka som köper något på en marknadsplats.
Ett litet barn som bär hjälm sitter i en barnvagn som ligger på golvet.
En flintskallig man i svart hatt klädd i svart skjorta med svarta skor på scen och spelar en röd gitarr på en konsert.
En man tar en bild med sin telefon.
Sett ur en låg vinkel, en man i en tank toppen spelar trummor.
Tre musiker uppträder tillsammans.
En stor gul skåpbil med en man bredvid på gatan.
En grupp på fyra vandrare i skogen.
En grupp människor i friluftsutrustning tittar på en karta.
Ett ungt barn på sjukhus dekorerar sin medicinska apparat för semestern.
En seriös man i en solbränd rock står utanför medan den snöar.
En liten pojke i en blå jacka förbereder sig för att skyffla snö.
Fyra vandrare går upp för trapporna på en liten kulle.
Man i blå skjorta sitter på sidan av vägen med en skottkärra av grönsaker
En tungset flicka i en randig klänning med glasögon håller hand med någon medan hon får någon form av medicinsk behandling.
En mor och hennes två barn sätter sig ner för att vila.
Två personer i gröna rockar och byxor, bär skyddsvästar och bär en stack orange kottar.
Ett par går upp för ett par trappor i snön.
Många hundar simmar och leker i en fontän i en allmän park.
Två män på byggnadsställningar fixar en fläck i en byggnad.
En man i en blå jacka kör en cykel laddad med en potatis typ grönsaker.
Kvinnor samtalar samtidigt som de sköter sina produkter på en marknad.
Två killar är i en soptunna och tre andra är i bakgrunden.
En kvinna som lutar huvudet på en mans axel.
Fyra personer i 30-årsåldern tar ett gruppfoto på en bar, någon flippar ur kameran.
Två personer i vita hattar tittar på en datorskärm.
En skäggig vit man i en mössa och gul jacka står bredvid ett fallet träd medan han tittar mot en annan man.
Skidåkaren i blått vänder och skapar ett dammmoln av snö bakom sig.
En kvinna i svart jacka tar en kopp kaffe.
Varmluftsballonger förbereds för användning.
En man med tatuering bakom örat spelar gitarr och sjunger in i en mikrofon.
Folk står på trottoaren bredvid vagnen och spår.
En halvcirkel av vuxna och barn sitter med en julgran i bakgrunden.
Två damer i vinterkläder som leker med en anka och snö.
En kvinna sjunger för en grupp människor som håller upp händerna.
Två asiatiska män jobbar med stålar.
Ett barn i en grön mössa sitter vid en båt kontroll.
En person går genom en snötäckt gata på natten.
En man i vit snöutrustning skyfflar snö.
En man i en gul lastbil som plöjer snö.
En kvinna bär håret ner och har inte huvudet täckt som de runt omkring henne.
Två män som arbetar utomhus på natten i snön.
En man som bär hatt håller en silverstolpe på en livlig trottoar.
Manliga och kvinnliga soldater lastar av julklappar från baksidan av en van.
Man och kvinna står bakom stor lastbil framför gult hus.
Två kvinnor kysser varandra vid en flod i en stad.
En grupp människor som försöker sig på skridskoåkning en solig dag.
En kvinna sover i baksätet på en bil.
En man skyfflar sina främre steg efter en snöstorm.
En man med röd skjorta lutar sig mot en motorcykel.
Hunden bär koppel i munnen rinner genom kärret.
Två personer går mot en kupolstruktur.
Två män i orange uniformer står framför ett tåg och gör lite arbete.
En kvinna och en ung pojke läste en bok tillsammans i ett vardagsrum.
En unge i gul skjorta brottas med en denim som bär barn på den vita soffan.
En man med grön skjorta tittar ner på en mobiltelefon.
Järnvägsarbetarna sätter fast ett band för att betjäna en bil på en lutning.
Folket marscherar genom gatan.
En man med blå skjorta vänder hamburgare på en utegrill.
En man håller en gitarr och talar i en monter mikrofon
En liten flicka med spetsiga flätor sitter i sanden på stranden.
Fyra män på en scen spelar olika instrument.
En man med skägg sitter på en klippa när han ser havet tvätta sig i land.
En polis mitt i en parad
Mannen i den svarta hatten har ryggen mot en teaterskylt.
Två äldre män pratar på trottoaren.
En man med blå och vit jacka, keps och ryggsäck, med fotografier.
Tre män diskuterar ett projekt längs sidan ett stort gult byggnadsfordon.
En brun valp som går genom snön.
En man och en hund går på gatan.
En tjej med svart hår och en brun tröja lagar mat på spisen och har ett stort leende i ansiktet.
En grupp människor som står i ett kök.
En tung man som bär hängslen sitter på en bänk bredvid ett stort ballongarrangemang.
En hund som springer genom ett fält mot en kamera.
En kvinna med blont hår njuter av solen i sin blommönster skjorta flip-flops.
En leende kvinna som sitter i en leende mans knä.
En person går uppför en snöig kulle med skidor på ryggen.
Ett litet barn som ler efter att ha begravts i sand.
Ett barn med röd hjälm, cowboyväst, randig skjorta, silvershorts och bruna byxor.
Ett par går genom regnet med sina barn som håller parasoller.
En man och hans far ser mycket roade ut som den yngre mannen i den blå skjortan och mästare hatt hålla upp en barbie docka.
En liten flicka leker klä upp sig.
En kvinna som står på gatan samtalar med en man på en lastbil.
Fem grundskolebarn kör en relätävling.
En flicka och pojke i blå tröjor passerar en stafettpinnen på ett spår möte i Asien.
En person driver en köttaffär.
Två unga pojkar håller ett gråtande spädbarn medan båda sitter i samma stol.
Två män i reflekterande västar går förbi en jättebild av en man i väst.
En utsikt nerför en smal europeisk kullerstensgata med flera bilar parkerade längs vägen.
En man kramar sitt barn på ett sjukhusrum.
En svept man som kommer ut från en mörk dörr och håller en skalle.
Två barn som kör ett relälopp.
Tre män i gula västar som gräver ett hål i jorden.
Tre män i en spricka på en gata.
En brun hund leker boll på en gård.
En kvinna som klättrar uppför ett berg.
Ett barn som bär en blå rock löper längs snön medan en liten hund följer efter.
Två män i tillfälliga kläder rör på sig krossade klossar av burkar.
Den nya lilla flickan somnade bredvid sina nytvättade och vikta kläder och filtar.
En publik sitter i en hörsal.
En gyrokock i vit jacka och keps som tittar på gyrokött.
En hane med röd hatt sitter på en stock i skogen.
En grupp människor tar en paus på sin vandringsresa.
En pojke i en röd tröja lutar sig mot en sten.
En ung pojke går igenom stora klippor i bergen.
En man står på en tunnelbana lutande mot en stolpe.
Här är en bild av asiatiska dansare som utför en ny dans framför sin klass och lärare.
Två personer hjälper en herre över vattnet.
En man läger utanför med ett tält och nödvändiga campingutrustning.
Två män filmar en äldre gentleman, medan en fjärde man tittar.
Ett litet barn som bär rosa sitter på en mörk matta.
En blond tjej som sträcker sig efter en korg leksaker.
En kvinna i röd t-shirt bär ett blont barn, medan en annan kvinna står i närheten i köket.
En pappa fixar en leksak åt sin dotter.
En kvinna med kort, mörkt hår står på golvet och läser en bok för en liten flicka klädd i vit klänning.
En mörkhårig kvinna kramar ett blont barn medan en kvinna i en fri skjorta klockor.
Tre personer i ett öppet utomhusområde har just landat från ett fallskärmsdropp.
En kvinna som går nerför en fullsatt gata
En man sitter ner pekar och tittar in i avståndet, det finns ölflaskor visas i bakgrunden också.
Flickan i blå klänning och hatt ler.
Ung barn gör sig redo att bowla en boll mot en nål medan du spelar bowling.
Sju personer går över en bro.
Två personer hoppar från ett plan och är på väg att släppa fallskärmen.
En basketmatch på college som spelas på konferensen "Stora tion".
En grupp människor pratar och står bredvid en busshållplats.
Tre klädda kvinnor går på en grusväg.
En asiatisk kvinna står vid en kassadisk och håller pengar i handen.
En tjej i rosa byxa som leker i marken.
En kvinna som shoppar knuffar sin barnvagn medan hon tittar igenom föremål på hyllan i gången.
Två män står nära en tung utrustning.
En grupp människor i formella kläder samlas i en kyrka.
En kvinna bakom ett glas ler och håller fredsskylten.
En ung pojke går över ett rör som rinner över vattnet.
Fyra barn som sitter ner två sitter på en vit duk.
Två lättklädda män sätter sig ner och njuter av en öl och mat utomhus.
Tre vänner ler för kameran eftersom de äter en intressant utländsk måltid.
Bredvid en grön fält, ung blond kvinna sitter utanför på en grå stammen applicera makeup på hennes ansikte.
En utförsåkningsåkare som bär en limegrön jacka och en vit hjälm.
En man och kvinna i formell klänning ler mot varandra när de dansar på en fest.
Fotbollsspelare i maroon jersey står bredvid domaren i svart
En fotbollsmatch i mitten av matchen, med en person i gult på väg att få bollen.
Tre fotbollsspelare står på ett fält.
Fotbollsspelare pausar ett spel eftersom en spelare i vit uniform skadas på fältet.
Den två mannen spelar softball.
En grupp människor i snön, en böjer sig över för att röra en snösko på hans fot.
Två unga kvinnor poserar stolt med snögubben de fullbordat.
En man i mörka kläder står bland några kugghjul.
En man springer mot en annan man som har fallit under en rodeotävling.
Idrottsmän på en fotbollsplan står runt varandra
En svart hund hoppar upp till en mans upplyfta hand.
Rodeo rider cowboy försöker hålla på en tjur i en arena omgiven av rodeo clowner.
Arbetstagare i orangea kostymer arbetar på en väg.
En man som sitter vid den offentliga tvättomaten och väntar på att hans kläder ska torka färdigt.
En korgie går på en tunn blå plattform.
En hona i violskjorta och svarta byxor är fokus för flera kameror.
En brun hund hoppar på bakbenen.
Åtta personer visas på bilden i snöutrustning som verkar vara skidåkning.
Två hundar står sida vid sida på gården.
Ett par som är väldigt glada över vad som pågår.
En man står vid en fruktvagn.
En kvinna i röd skjorta står ensam i en terminal, med tre bagagelappar.
Tre kvinnor klädda i grönt och shamprocks.
En medelålders man med en knapp upp skjorta läser en bok om hundar för ett litet barn som sitter i hans knä.
En mor, som lär sin lilla flicka.
Två flickor försöker korsa gatan i en fullsatt asiatisk stad.
En man står framför en spegel.
En liten brunhårig pojke med röd skjorta och blå jeans bär en grön lastbil.
Två unga pojkar leker med två små flickor.
En ung pojke i röd skjorta spelar i ett träd.
Tre tonåringar dansar en kväll på gatan.
En man sover på en parkbänk.
En husfest full av unga människor.
En man kastar något i en flod i staden.
Skidåkare i orange jacka, stående på toppen av en kulle
En ung person spelar gitarr, bakom dem står en mycket ljus lampa.
En man i väst står på en lugn gata.
Tre barn klädda i vinterkläder går genom skogen medan de driver med lasten.
En byggnadsarbetare i en röd hatt tittar på en maskin.
Många människor går nerför en gata omgiven av gamla byggnader.
Kvinnan inlindad i filt sitter på bänken och läser i parken.
En röd hattad man styr en röd maskin för att rensa ut vägen, med blå himmel och grön stress bakom sig.
En bebis i gul skjorta ler.
Arbetare förbereder mat för människor att äta.
Någon i en röd skjorta som staplar många djurhudar.
Fyra äldre män spelar musikinstrument i en park vid en vägg i traditionell kostym.
En äldre man väntar på en tur på en landsväg.
Två äldre män står framför en butik av olika slag.
En man i förkläde använder butiksutrustning.
En grupp fotgängare går nerför en stadsgata.
En kvinna med en vit hästdräkt och hjälm tycker om att umgås med vänner.
Mannen i kostym med rosa skjorta och randig slips ger ett tal medan andra skrattar.
En elektriker som arbetar med ljus, möjligen luftkonditioneringskanaler i en kontorsbyggnad.
En man vilar på vägkanten med sin kamel.
Två personer som fiskar med en båt på bryggan.
Någon klädd i en grå topp ser på när skålen rullar ner längs fil åtta på den färgglada bowling gränden.
En man rider en häst i en parad.
En grupp människor stirrar åt samma håll och en kvinna sitter på en annan kvinnas axlar för att ta en bild.
Ett barn ler när hon klättrar.
En man i vit mössa, stående i ett fält med en fladdermus, på väg att svinga mot en boll.
En apa klättrar över ledningar ovanför en gata.
En man i snön på en ramp som arbetar på en isskulptur.
En professor undervisar en stor grupp studenter.
Tre unga män tar en bild på två flickor i en bar med en kameratelefon.
Ung flicka som gör sig redo att klättra.
Man i tung svart rock röker cigarr står nära kvinna i brun jacka med ett papper i handen
En hund som går längs en snödriva.
Det finns många människor som går runt och tittar på saker i det röda rummet
En man i kostym står bredvid en stor målning omgiven av en stor guldram.
En grupp människor på en buss eller en tågbil.
Två personer som bär snöskor hoppar upp i luften för att posera för ett foto.
En man i orange och grå jacka som hoppar i skidor.
Två personer sitter på en brygga med en solnedgång i bakgrunden.
En man och en hund på en parkbänk i förgrunden, med en grupp promenader människor på avstånd.
Två små barn som bär vinterkläder skyfflar snö.
En man sitter i en stor blå båt och tittar på smutsigt vatten.
En blond man med ryggsäck står bredvid en damm.
En pojke drar en liten pojke i en röd släde genom snön.
Folk går och äter framför ett hotell.
En grupp människor som försöker dra en traktor.
En häst som tar en cowboy i rodeo
En kvinna i röd jacka, med en hatt och halsduk på huvudet, säljer sina kläder på trottoaren.
Två män rider på en tunnelbana medan de läser böcker utan byxor.
En flicka i vit stickad hatt och vinterutrustning gnuggar tungan över tandställningen.
En man väntar på att få en drink från en flygvärdinna.
En man och en kvinna diskuterar nåt över drinkar på en bar.
En man pratar med män vid ett bord.
Rodeofolk går ut genom en grind med en kvinna och en pojke som följer efter dem.
En man skateboardar i en stad.
Ett barn knuffar eller sparkar en fågel med foten.
Ett gammalt par spelar musikinstrument i ett gathörn.
En skäggig man läser medan han sitter på en vägg i en park.
Två herrar står utanför en Smoothies &amp; Bubble Tea försäljare.
Två stora koner är utanför, på gatan, framför en stor byggnad.
Ett par pojkar är i ett gym med delvis monterade cyklar.
Två män på motorcyklar, den ena med silverhjälm och den andra med svart hjälm, ridande i en stad, med en pojke med en vit långärmad skjorta på, närmar sig en av motorcyklarna.
Elever, och deras lärare i ett klassrum går igenom material.
En hund springer på ett fält med munnen öppen.
En brandman har visat sig försöka klättra in i några spillror.
Människor som samlas längst fram i templet innan de går för att meditera.
En man i vit skjorta närmar sig en mås.
Tre kvinnor är utanför och en av kvinnorna ler.
En man erbjuder prov på mat.
En kvinna som går ut medan en gentleman rider på en motorcykel i närheten.
Två män med nyanser som pratar på balkongen.
En kvinna läser en bok för två små barn, en som dricker ur en kopp.
En man i gul skjorta leker med sin svarta pudel.
En man i en ljusblå skjorta och khaki shorts som håller en vattenflaska går nerför stigen mellan två branta grottväggar.
En flicka klädd som en fjäril.
En skateboardåkare flyger genom luften medan två personer observerar från en lång utsiktsplats.
En wakeboardare utför ett trick på en räls.
Framtiden för snowboard på sommaren med all den höjd och spänning du kan önska dig.
En ung hane gör ett cykeltrick på en bro på kvällen.
En grupp människor hoppar iväg på en gata
En extrem cyklist skär ett hörn i skogen.
Två unga flickor i ett kök som bär förkläden över pyjamasen hälsar en man i en olivgrön skjorta.
Det här är en kvinna som spelar sin flöjt med noter framför sig.
En man klädd i grönt med ansiktet täckt av en bandanna arbetar utomhus med tunga maskiner.
En arbetare vilar foten på baksidan av en husvagn.
En man som bär en tågledares uniform stående inuti ett gammalt tåg eller vagnsvagn.
Kvinnan med en röd hatt skridskor och går sin hund.
Åskådare tittar på hästar och deras ryttare på en inhägnad stig med en damm bakom stigen.
Jag unga flicka blåser en bubbla med tuggummi.
En liten asiatisk pojke bär gröna pärlor och håller i en grön Saint Patrick's Day ballong.
En sky-vy av män som gräver hål genom betong.
Två män står vid en lastbil och bitar av trädstammar.
Skäggig gammal man har diskussioner på vagn.
En grupp afrikanska barn klädda i olämpliga kläder sjunger och spelar instrument.
Två personer går på en gata med karga träd.
Närbild på sidan av en gammal kvinnas ansikte med överdimensionerade solblockerande glasögon, grått hår och ett guldörhänge.
En ung, asiatisk man ses spela gitarr.
En man som bär en långärmad, blå rutig skjorta och bruna byxor knäböjer bredvid en hjulvagn i ett garage.
En man håller fast ett blöjat, blåskjortat spädbarn på knät.
En man och en kvinna pratar med varandra över ett skrivbord.
En byggarbetsplats sliter sönder en vägg med graffiti.
En brun hund jagar en röd frisbee över ett gräsfält.
Två barn sitter vid ett skrivbord.
En grupp människor sitter vid ett bord och äter tillsammans, de är i en fin restaurang.
Bilen lämnade ett stort rökmoln.
En Volkswagenbil kör genom ett ökenlandskap mitt i bergen.
En kvinna som lagar middag hemma.
En grupp människor lyssnar på en man som står på ett podi.
Fyra personer vaknar i snön utanför.
En man klädd i vinterkläder som hugger ner ett träd i ett snöfyllt fält.
En grupp löpare som avslutar ett lopp.
Tjejen springer i ett maraton, bär en svart skjorta med en vit tank topp, med nummer 44 på.
En blond pojke i randig skjorta som ska sparka en rosa fotboll.
Människor som står framför en grå byggnad med en skylt som lyder 'Tickets Tillgänglig Här'.
En kvinna med tårfläckat ansikte på ett piano.
En man som använder skidutrustning hoppar genom luften nära en tegelbyggnad och blå skyddsräcken.
En brun och vit hund hoppar, håller en flexibel Frisbee.
Ett lag i röda och svarta uniformer står på varandras axlar medan folkmassor pressar in dem.
En kvinna och en man står utanför en affär.
Ett band spelar ute på en stengång.
Många människor samlas runt gatan och tittar på två gatuartister.
Fyra kvinnor samlas i traditionella klänningar och tittar på ett evenemang.
En man som rider på en häst och tävlar om att bli nummer 1.
En man tvättar eller dör kläder i en primitiv miljö.
Män som arbetar i smutsiga förhållanden med rött tyg.
En kvinna som lagar mat i ett förkläde ler mot kameran med två andra kockar i bakgrunden.
Två personer klädda i svart vända bort från kameran med skallben på sin jacka respektive ryggsäck.
En man har en mikrofon, medan ett par dansar i närheten.
En svart hund som leker med en grön leksak.
I folkmassan finns en kvinna i en röd rock längst ner i trappan.
En grupp unga musiker.
Ett band som inkluderar en Upright Bass Player spelar i ett tält framför kanadensiska flaggor.
Ett band gör sig redo att spela.
Nio kvinnliga dansare bär tutus och använder "Guitar Hero"-gitarrer som rekvisita på scenen.
Män som gör sig redo för SXSWO att gå live i sändning
En man i blå skjorta och svart huva tittar på en annan man, i en blå skjorta, gör något med elektronisk utrustning.
En man som bär vinterjacka tar en bild.
En person sätter sig i en bil parkerad framför Swan Restaurant i snön.
En ung orientalisk pojke som håller i en trumpet som pekar åt höger.
En svarthårig kvinnlig gitarrist och en manlig trummis spelar i ett stort tält.
En man spelar mini-guld på SportsCenter set medan två andra observera.
En pojke hoppar på en stor hög löv medan en grupp barn och en kvinna tittar.
En man petar på en eld med en pinne medan han ler.
En kvinna och två små flickor sitter på en betongbänk med händerna på läpparna.
Två arbetare sopar trottoaren utanför sin lilla affär.
En gränd öppen för ett par människor som går förbi
En kvinna bläddrar igenom några prydnader.
Ung man i kamouflagebyxor bär en stor metalllåda som går längs trottoaren.
Två turister fotograferar en landsbygd och ruiner
En afroamerikansk man som står med ett blått träkort med två hjul på en sandstrand.
En man ligger ner i gräset.
En man i kostym pratar på en directtern.
Tre män pratar på en entreprenörsmässa.
Två män står och pratar med varandra, en av dem bär en skjorta som säger "sommarskola".
Två män som tittar på tre kvinnor som tittar på en produkt.
Tre personer sitter vid ett litet bord nära en skärm med orden "DEMOS, The Business of Care".
Tre personer sitter vid ett bord framför en folkmassa.
Kvinnor som står på podiet och pratar i en mikrofon.
En stor grupp samlas för en bankett.
Folk i kostym står vid ett bord med en röd duk.
Pojken i shorts badar med slang på gatan.
En äldre kvinna som bär en grön jacka och en röd hatt håller sin svarta axelväska när hon tittar på avstånd.
Personer som äter en McDonalds-måltid längs gatan.
En äldre kvinna i glasögon och en vit och svart skjorta som arbetar med färger.
Två män går, en med hund och en bajsscooper.
En kvinna som bär en blå jacka står utanför bredvid en cykel.
Folk står i en park bakom en prydnadsbåt.
Ett litet barn använder en slipmaskin när de bär skyddsglasögon.
En lärare som hjälper en liten flicka med en maskin.
En man med huvudet nära en laptop som trycker på en knapp.
En kvinna sätter ihop ett träföremål.
En ung flicka bär gula shorts och en vit tank topp med hjälp av en käppstång för att fiska vid en liten damm.
En hund fångar svart Frisbee.
En grupp människor framför ett skyltfönster klädda i vinterkläder på kvällen.
Två äldre människor tar en promenad längs en trädkantad stig.
En orange lastbil ses som food trucks rad upp på en gata.
En man som ristar upp kött till en måltid.
En äldre dam med röda skor, rosa halsduk, grå hatt, och hålla en väska, föra ett samtal med en äldre man med röda byxor, grön rock, och en grön hatt.
En man utanför en mobil lunchbil.
En gammal afrikan med en cigarett i munnen som sitter med en maskin framför sig.
En grupp elever som arbetar tillsammans i ett klassrum.
Ett mycket litet barn gör ett surande ansikte på en äldre hane i en skinnjacka.
En man och kvinnor är på en buss.
En ung flicka sitter i fosterställning i smärta.
En asiatisk man med långt vitt skägg som stirrar rakt fram.
En blond kvinna i högtrycksskjorta som höjer handen och ler.
En stor publik är närvarande vid ett evenemang och tar bilder.
Folk ser på ett monument där en hastighet ges.
En blond man sjunger och spelar gitarr.
En man håller upp en liten klistermärke som säger "Jag är en fotograf, inte en terrorist" medan står bland en stor grupp demonstranter.
En dansare som uppträder med en hulahoop, med domare i bakgrunden.
En ung kvinna är med i en gymnastiktävling.
En ballerina framför en jury av domare.
Hantverkaren sitter utanför och arbetar med sin trampmaskin för att fläta rep.
En kvinna ler och håller upp en Spindelmanskjorta.
En man och en kvinna sitter på golvet och arbetar med pysselföremål.
En grupp små barn i en by utan asfalterade vägar.
En stor skara människor som sitter i läktarna och tittar på en fotbollsmatch.
En man som bär halmhatt hamrar något.
En grupp män och kvinnor som tittar på konst i en konstutställning.
Ett litet barn bär några roliga glasögon som är alldeles för stora för hans ansikte.
Ett par människor på ett museum tittar i presentbutiken, potentiellt kommer att köpa något.
Killen på cykel med ögonen tysk Shepard hund.
En husky-hund sniffar en hästs axel medan hundens ägare klappar de två bruna hästarna.
En man som bär en blå jacka visar glatt sin produkt.
En kvinna med glasögon kammar igenom håret med fingrarna när hon skriver i en anteckningsbok med en penna.
En ung flicka som skriver med en lila penna.
En kvinna hukar sig ner för att nå en hink full av döda och skinnade kycklingar.
En grupp människor sitter under paraplyer på stranden.
En person, klädd i en röd jacka, åker skidor nerför ett snötäckt berg.
Byggarbetare sätter ihop ett vitt tak.
En sjuksköterska övervakar ett litet barn som verkar vara post-op.
En person som bär grön skjorta hoppar på sängen.
Två kvinnor, en äldre och en yngre, tycks vara ombord på kollektivtrafiken.
Två unga pojkar äter sin lunch utanför på cementtrappor.
En kvinna sitter i en stol och ler medan hon håller ett sovande barn.
En kille som får pengar från en bankomat.
En publik som står i grupper på cementområdet mittemot parkeringen och bygger i bakgrunden.
Den svarta hunden retreiverade den vita leksaken i vattnet.
En kvinna i svart uniform trycker ner en gul mopphink i korridoren.
En sittande man som spelar fiol.
Tre killar bär pyjamas, två sveper golvet medan de andra tittar i ett klassrum.
Två kvinnor de båda bär en mörkblå uniform
En person som bär en blå och vit rock cyklar nerför gatan.
En man klädd i rött spelar gitarr på en gata.
En liten flicka i rosa klänning lägger huvudet på en kvinnas knä och suger i tummen.
Två män står bredvid ett matstånd.
Flickan paddlar en rostig kanot i vattnet.
En man stickar äger några maskiner.
En man tar en svandykning från en klippa medan andra tittar på.
En man i vit skjorta jobbar vid ett bord.
En vagnsbil passerar genom en stad.
Barn äter popcorn medan de sitter på bönsäckar.
En arbetare tittar på sin laptop som sitter vid hennes skrivbord.
Hunden hoppar över baren.
En löpare är på väg att springa under bron i höst.
En man som sitter inne och tittar på fönsterputsaren utanför.
Två killar på en soffa, den ena tittar upp den andra tittar bort med en kopp i handen.
Den bruna hunden springer i vattnet och slickar näsan.
En buss öppnar dörren för att släppa av och av folk.
Två barn sitter vid ett skrivbord medan en annan sitter i fönsterbrädan.
En bild av en liten pojke på en trottoar som tittar på en duva.
En stor kvinna i en blå jacka ser irriterad ut.
En man och en kvinna sitter på en buss, men inte tillsammans.
Ett litet barn som bankar en plasthammare mot en metallkruka.
En kvinna som bär en fanny pack tar ett foto av en röd bil.
En häst eller mula drar en man i en kärra nerför en asfalterad väg.
Tre cowboys rider sina hästar bredvid ett staket, i en torr gräsmark.
En simmare i en blå baddräkt ler för ett foto.
Två män hoppar över en stor blå vattensamling.
En basketmatch innan den börjar.
En grupp människor sitter på en basketarena och tittar på ett lag som bär blå och gula tröjor som värms upp.
En ung man spelar piano och sjunger på en konsert.
En man i grå t-shirt och svarta shorts som håller vad som verkar vara hans son.
Ett barn sover på en filt.
Sport lagmedlemmar öva och koppla av på en basketplan.
Kvinnliga basketspelare värms upp innan ett spel.
En grupp människor, mestadels tonåringar, arbetar på en trottoar, gräver och städar upp vinstockar.
Två kvinnor som håller spadar står på en liten bergssluttning.
Ett litet barn i vinterkläder hoppar i ett snöigt och trädbevuxen område.
Mannen står på gatan och håller en skylt
En man rakar ansiktet medan han tittar i spegeln med rakkräm som täcker ansiktet.
En vuxen kvinna och en ung pojke går genom en stad på kvällen.
Gymnast ligger på golvet med ett ben pekat upp i taket.
Brun hund som hukar sig i gräset och tittar upp
En man i en knapp upp skjorta spelar xylofon.
Unga flicka tar låg hängande telefon medan en man går iväg.
En grupp fotbollsspelare på ett fält, det ena laget bär svarta och blå uniformer, det andra rött och vitt.
Människor i vackert blått vatten surfar en fin våg.
En flicka som bär en rosa skateboardhjälm rider i en skateboardskål.
Ett olyckligt barn som ser ut att ligga i gräset i en park.
Tre personer, som var och en bär ett par röda snöskor, slappnar av i snön.
Två bruna och vita hundar i gräset nära en stenstruktur.
Ett barn med blont hår tittar på ett urval av kakor och brownies.
Hunden är framför några buskar.
En stor grupp män lyssnar på en man med glasögon som sitter vid ett bord med ett konstigt mönster.
På det här fotot ler en kvinna i telefonen.
En man i blå rock och jeans äter en korv.
En tjur laddar en matador i rodeo, medan tre andra män tittar på djuret.
En tjurryttare är i luften och ramlar av tjuren som är i bakfoten.
Två människor ler medan de slädar nerför en snötäckt stig kantad av tallar.
Fem män i tung vinterklädsel som rider nerför en snöig kulle.
En vandrare använder metallstavar för att vandra uppför ett snöigt berg.
Ett olyckligt barn med slutna ögon rör vid någons byxor.
Tre barn är vid en vattenväg bakom ett hus.
Ett litet barn i en vit huva jacka håller i sig mot väggen.
Åtta orientaliska tonåringar i röda skjortor sitter på betongblekar.
Ett litet barn som bär blå jeans och en vit skjorta ligger på marken längs sidoutskurna pappersträd och en sol.
Eleverna är i ett klassrum och läser något från en tidning.
Det finns flera asiatiska barn som sitter korsbenta på ett betonggolv.
Två tjejer äter en måltid tillsammans.
En ung pojke tar en tupplur under en kartong som lyder "Connie Facial Tissues".
Asiatiska skolbarn presenterar ett gruppprojekt tillsammans.
En pojke tittar på ett märkligt lila föremål i sina vänners hår.
Fyra barn som spelar basket i ett gym.
En mörkhårig flicka som håller i ena handen och visar fredsskylten med den andra handen.
Fyra studenter sitter på golvet vid en modellvulkan.
En grupp asiatiska elever spelar London Bridges medan en annan elev ligger på marken.
Två unga elever som delar med sig av sina uppgifter inför klassen.
Två asiatiska elever försöker pussla ihop något.
Ett musikband som spelar musik.
En grupp unga människor som alla bär röda skjortor och alla bär väskor eller plånböcker.
Folk går in i en väldigt lång, gammal byggnad.
Asiatiska gymnasieungdomar gör en gruppaktivitet i en cirkel.
Asiatiska studenter undersöker pappersark medan de står i kö.
En ung asiatisk flicka har en uppstoppad kattleksak i ett klassrum.
Tre ungdomar står i ett trångt rum.
Två flickor sitter vid ett bord med en grön markering som står på dess ände.
Eleverna läser sina svar i klassrummet
En grupp unga flickor sitter på en buss med de flesta tittar ut genom fönstret medan man tittar på kameran och ler.
En klass elever som alla gör olika handlingar.
Barn som leker i ett gym med ett dukväggsöverdrag på en vägg.
Fyra asiatiska barn sitter på golvet i ett klassrum.
Två flickor skrattar leende när de sveper in ljust färgade snören i varandras hår.
En kort man håller tal.
En tjej i blå klänning spelar på en lekplats.
En okänd solider i grönt pekar på sin högra visar en annan man något
En grupp människor som bär orange och svart spelar olika typer av trummor som andra tittar på.
En grupp välklädda ungdomar står framför en församling.
Två män står i snön, en tittar på kameran, den andra läser ett papper med en skylt.
Två män åker skidor och den till höger skrattar.
En man i svartvit baddräkt, ser ut som han hänger i luften, gör sig redo att hoppa i en bakgård pool.
Både män och kvinnor är vagt klädda, med sina armar sammanflätade mellan varandra.
En kvinna dansar i löv, medan åskådare sitter eller står på gräset.
En man står ovanpå ett byggnadsfordon.
Barn leker på trottoaren nära en adobe byggnad.
En man på kryckor läser tidningen.
En baby spelar schack som en katt tittar på.
En man som bär växter och örter längs en tågbana.
Ett ungt, blont barn tittar ut genom en glasdörr.
En ung man som står under ett Playboy-tecken.
En bonde tar sina apelsiner till marknaden för att sälja.
Många cyklar är parkerade bredvid varandra.
Skolbarn klädda i uniformer ser sig omkring i sin omgivning i klassrummet.
Barnet sover medan han äter.
En massa människor klämmer genom flygplatsen.
En man och barn som tar emot saker från en kvinna.
En lång man klädd i långärmad skjorta, byxor och långa stövlar sveper på en gård.
Två kvinnor tittar på bröd på ett bord.
Två kvinnor i kjol står bredvid en byggnad av sten.
En ambulans är nära en tall.
En man spelar gitarr och två kvinnor i korthet, vita klänningar står bredvid honom.
En mor som gärna drar sitt barn i snön med en släde.
En man som står i brun jacka och skyfflar bort snön från vandringsvägen
Två manliga barn städar upp löv på en parkeringsplats.
En vuxen dam som bär en tanktopp och en kjol ställer disk i diskmaskinen.
En man med skjortärmarna rullade ihop gester medan han talade.
En skidåkare i röd snödräkt och vit hatt håller i en skidstolpe medan han står i snön.
En man serverar mat till en pojke.
En man som bär rock och floppy hatt trycker en blå kundvagn full av väskor.
En man som bär hatt är bakom ratten på en vit propanbil.
Ett snötäckt landskap med ljusa armaturer och ett rött staket.
Människor vandrar genom ett isigt, kuperat landskap.
Tre män, klädda i regnkläder, står på en båts brygga och förbereder sig för att rena fisken.
Hundägaren försöker hämta frisbeen från sitt husdjur.
En grupp män och kvinnor som äter och dricker.
En man och en kvinna står på trapphuset
En grupp barn som står runt en staty i en lobby.
Barn sitter på en vägg inuti en kyrkogård.
En man tar en bild medan en annan tittar på i en utländsk butik.
En kvinnlig sångare uppträder på scenen.
En man sitter vid ett bord och pekar medan två kvinnor tittar på honom.
En flicka som går nerför trottoaren på natten
Tre personer står vid en strandlinje och har ett stort nät.
Folk sitter runt ett bord med menyer och vinglas.
En person som bär en tonårings kläder och en ryggsäck ligger med ansiktet nedåt på en vadderad bänk.
En man i grå skjorta känner sitt skägg.
Män och kvinnor som står på en bräda och sätter upp sidospår.
En man sitter på en cykel lastad med lådor.
En man som spelar gitarr och sjunger med en annan man
En kvinna tittar på bilder i ett fotoalbum.
Två unga män brottas med varandra mitt i ett fält.
En skateboardåkare gör ett trick i luften.
Flera män och kvinnor klädda i orange västar går på en snötäckt väg på vintern.
Två kvinnor som sitter på golvet och gör filtar.
En man i röd skjorta betjänas av en arbetande gammal kvinna i en affär.
Tre män väger fisk när de kommer av båten på en skala vid kusten.
Underhålls- eller byggnadsarbetare på en arbetsplats på en livlig stadsgata
Äldre kvinnor i en blå tröja som spelar piano vid fönstret.
En äldre man som tippar på hatten medan han står i en grupp människor.
En grupp proffs som sitter runt ett bord.
En man ställer upp för en väntande smet när de spelar på en parkeringsplats.
En man står utanför ett hus med en snöskyffel.
En man i svart cape vänder sig mot en ung pojke i träningsoverall.
Ett område är täckt av snö.
En man och kvinna står framför en stor röd modern staty.
Pottery kan avnjutas av även de mycket unga i hjärtat.
Barn blir besprutade av en vattenspridare.
Mannen knäböjer på biltaket och hjälper till att lossa ved.
En ung flicka i en lång rosa blommig klänning och matchande headscarf går ut och bär två stora, fyllda, vita tygpåsar, en i varje hand.
En riktig cowboy, den här mannen håller i sig under ett spännande rodeo ögonblick.
I en parkscen hoppar en man över ett föremål på en skateboard medan en annan man knäböjer med en kamera för att ta ett foto av hoppet.
En ung kvinna som bär polotröja och svart jacka ler för en bild.
En kvinna poserar bredvid en bur full av uppstoppade hajar med tecknade serier målade på väggen bakom henne.
Två killar övar på handslag.
Lilla flicka med brun snöjacka och lila snö byxor leker i snön med en röd spade.
En skjortlös man håller i en ansiktsmask.
En äldre man plockar upp bitar av trasiga barbiedockor.
I Ikeaaffären sitter en man på en stol.
En grupp damer som går längs en trottoar bredvid en blå och vit vägg.
Två pojkar i stora bubblor på vattnet.
2 spädbarn, 1 i varm rosa jacka och andra i rosa och blå blomjacka kramas i snön.
Går hem en kall vinterdag.
En grupp människor som har bråttom att börja arbeta.
Två män i clownmakeup gör en musikskit på scen.
En kvinna sjunger på en scen medan en man i clownmakeup spelar gitarr.
Ett barn sover och suger på fingret.
Fyra bandmedlemmar spelar på en röd scen framför ett stort hjärta.
Tre musiker uppträder på en scen upplyst med rött ljus.
En kvinna med ryggsäck och en akvagrön skjorta med handen på huvudet och hennes hår drog upp tittar över några kullar.
Ett barn leker i snön med en grön spade.
En man i svart och vit randig skjorta sover på en betongbänk.
Två små flickor cyklar.
En kvinna i svart tank topp och shorts går längs sidovatten medan hon lyssnar på sina hörlurar.
En svartklädd man spelar munspel.
En man som undersöker vad som verkar vara mat i ett kök.
En baseballspelare förbereder sig för att svinga slagträet på en boll.
En bagare klädd i vitt med en hårnät fungerar med deg med hjälp av en lång stolpe.
Två kvinnor som sitter på ett trapphus i en mestadels vit kakelbyggnad.
Man i mörka kläder när han står framför en upplyst julgran i skuggorna.
En man som står framför en ugn med bröd i.
En man, som svingar en kniv, tittar på mat på en rotisserie medan andra ser på.
Ett mycket litet barn bär en vit dräkt runt huvudet.
En asiatisk man sitter ner med ledningar som kommer ner med en resväska bredvid honom med bilder på kvinnor på.
Två män går bort från en bänk.
En kvinna i en svart tröja häller flytande tvättmedel i en tvättmaskin.
Svart hund som springer genom ett gräsområde.
En kvinna som just avslutat sin dansföreställning3.
En brunhårig man som sjunger medan han spelar gitarr.
En kvinnlig gymnast är upp och ner med benen i delad position.
Två poliser cyklar på gatan.
Två unga flickor med långt hår som ler med rosiga kinder, en med röd skjorta, en med vit skjorta medan de gömmer sig bakom en vägg.
Två personer bär sina väskor på en obesegrad väg.
En pojke går i snön med sin hund och håller sin snowboard medan en äldre man, förmodligen hans far, följer efter i bakgrunden.
En tjej med vit och röd makeup som håller i ett rött paraply.
En grupp på 4 personer går längs en stig.
Tre män i en liten båt sänks ner mot vattnet.
Barn och vuxna bär vinterklädsel ridande cyklar nerför gatan.
Två personer sitter på en sten i en stads park.
En brun hund försöker fånga en flygande skiva men missade den.
En man som går runt hörnet av en röd byggnad.
En man med byxor är på en bergsvägg.
Två kvinnor äter mat tillsammans.
En man i orange jacka tittar på stenar staplade i kolumner.
Athlete kastar ett spjut på ett spår och fält händelse.
En fårhund håller på att granskas av domare vid en hundutställning.
En publik tittar som fem hundar bedöms på en hund show.
En man som bär en blå skjorta står på en orange stege för att fixa ett ljus
En person i blå leggings njuter av skridskoåkning.
En kvinna på en buss som inte ser så glad ut och bussen verkar full.
Många människor på en hundutställning på en stadion.
Människor i linje med sina skidor på en skidort.
Två män klättrar på en trä byggnadsställning.
Tre personer i rockar som går längs en snösträckt stig på ett berg.
Tre personer med sina schäfer går på en grön gräs.
Ett barn stirrar utåt bakom en järnlaterad barriär.
En kvinna som ler bär en unik huvudprydnad.
Person klädd i mörka kläder gör en vända in i snön längs sidan av vägen.
En brun hund visar tänderna.
En beagle och ett ungt blond barn som bär nummer 96 på ett evenemang.
Herrarna med en snobbig jacka målar det omgivande landskapet vackert.
En man och en kvinna i färggranna kostymer utför en dans på natten.
En ung flicka och en tysk shepard på en strand.
En mor, hennes barn och deras hund är på stranden och ser ut som om de är på semester.
Ett asiatiskt par står vid en fantasiaffisch.
Tre personer i kroppsdräkter ligger på marken och verkar skrika.
En man lägger armen runt sin flickvän på en konferens.
En grupp människor i ett rum som pratar och sitter i stolar.
Folk serverar sig själva mat på en buffé på natten.
En man i vit jacka håller en pojke, som också bär en vit skjorta, i sitt knä.
Två tjejer spelar en sport.
En äldre man målar en landskapsbild som är på en staffl utomhus.
Mannen sitter på en sten med ryggsäck och en halsduk runt sin nästa ser ut att vara ledsen.
En man i en grön rutig skjorta som uppträder lite karaoke med gitarr framför en liten publik.
En man som pratar med en grupp människor.
En man och en kvinna, båda håller paket, pratar med två sittande män i ett väl upplyst lobbyområde.
Talare i ett rum fullt av folk som sitter i stolar.
En man i vit skjorta och jeans som använder en motorsåg för att hugga ner ett träd
Ett barn med vit jacka stående i snö.
Två personer tar sin båt ut i havet.
Ett par kyssar framför ett stort ishjärta.
En sju person som kallas soljägare leker utomhus med en skylt som ber om donationer.
En person i röd och guldklädd dräkt står bakom en man i svart.
Folk i en buss som är på väg till 84 Peterson.
En man och en kvinna arbetar med ett verktyg på en logg.
En gammal kvinna i huvudbonaden tillsluter marken på ett fält med hjälp av en hake.
Ett barn tittar på en ödla i ett annat barns hand.
Medan han sjunger in i mikrofonen spelar mannen i den svarta skjortan en akustisk gitarr.
Två män, en kanna och en umpire, är utanför och spelar baseball.
En manlig snowboardåkare som bär orange och blått stående ovanpå ett blått bord på en skidort.
En grupp människor samlas i en park under vintern.
En kvinna vilar på trottoarkanten på en stadsgata medan hon pratar på sin mobiltelefon.
En man går på en trottoar som håller på att byggas.
Två unga pojkar spelar spelet "Twister" och har placerat sina händer och fötter på blå och gröna fläckar.
Flera människor kör ett lopp.
Mannen med blå hjälm rider på en Polaris.
En ung flicka som gör hantverk, medan några människor står och tittar på.
En kvinna med svart bälte gör någon form av kampsport.
En kvinna som sitter vid en snurrande vävstol.
En ung indisk pojke blåser bubblor med en klassisk bubbelblåsare.
En ensam fiskare är på sin båt och kollar nätet.
En kvinna från Indien som stod och tillverkade garn.
Folk samlades runt en olivhandlare på en bondemarknad.
En man i mörkgrön jacka liftar en svart häst till en svart stolpe.
Berget klättrar nerför sidan av en stenig klippa.
Ett affärsevenemang äger rum med en attraktiv blond kvinna som ler mot kameran med sin telefon i handen.
Folk går nerför en gata med en gul moped i förgrunden.
En skridskoåkare håller den koreanska flaggan medan han vinkar till fansen.
En kvinna med nummer 145 kör ett lopp.
En spansk man som bär svart håller handen på en dansande kvinna som dansar.
Fyra barn sitter i ett pastellfärgat klassrum.
Detta är bilden av sex asiatiska barn med tamburiner.
Ett barn i denimjacka spelar hus.
En ung flicka som står framför en rad gula stolar.
Fyra kvinnor interagerar på en konferens.
En kvinna håller i nacken och tittar på något.
En mörkhårig kvinna på mobilen har en liten flicka i rosa klänning.
En hemlös man ligger på marken med sina grejer strödda runt.
Joggare i ett lopp en kall dag.
En stor grupp människor i ett rum, ler och skrattar.
En grupp kvinnor står och tittar åt samma håll.
Folk klappar händerna efter talet.
En kvinna i svart lägger armen om en annan kvinna medan de fotograferas.
En maratonlöpare som antingen startar eller passerar genom en vägspärr vid en insamlingsmaraton.
En skara människor förbereder sig för ett maraton.
Runners fotograferas som åskådare titta på och ta bilder av en Run för Haiti.
Runners tävlar i ett maraton.
En kvinna bär skridskor och det finns grupper av människor i bakgrunden.
En man kastar en lök i luften i köket.
En man och en kvinna går nerför gatan en kylig morgon.
Flera små flickor är på en bordsmålning.
Ett par dansar medan andra tittar på en konsert i ett bandställ.
Folk springer i ett maraton.
En tjej i hatt sitter på en strand medan hon pratar på mobilen.
Maskinen gräver ett stort hål på marken.
Marathonlöpare är på väg genom en park en kall vinterdag.
Runners tävlar en kall dag i stan.
En man som går barfota ser på över en klippa när solen är precis ovanför horisonten.
En skäggig man utan t-shirt fixar sin cykel.
Folk står i kö vid en vit bordsduksklädd buffé och serverar sig själva mat.
Två små barn går iväg på ett fält.
En grupp unga och äldre människor samlas runt om och håller i sig ett fridsamt täcke.
Ett stycke väggkonst som innehåller ett träd
En liten flicka i en vit tröja med prickar leker med ett träspårat tågsätt.
En liten flicka som kollar hennes kläder.
Två mörkhåriga män i orange skjorta som lutar sig mot ett skrivbord bredvid en man i uniform.
Ett lyckligt barn sitter i knät på en kvinna som bär en grön skjorta.
En person i orange skjorta ligger på marken medan andra står runt henne och ler.
Barn uppträder på en scen med tält i bakgrunden.
Det finns tre pojkar på scenen med podier framför dem, de förbereder sig för ett tal.
Två pojkscouter i jeans uppträder på en scen med tält.
Fem killar sitter på en scen framför två gröna tält bakom en scout av Amerika banner.
Pojkscouter på en scen med mikrofon
En ung pojkscout sitter i en campingstol framför ett grönt tält, inomhus.
En man går i en klargul jacka.
En ung orientalisk flicka i en rosa och grå randig skjorta nafsar på en jordgubb när hon tittar på henne rätt på något bakom kameran.
Två personer har picknick vid en sjö.
En man i orange väst står bredvid en gul kanot.
En grupp pojkscouter som ger en demonstration.
En grupp scouter står i kö.
Två tonårspojkar i pojkscoutuniformer.
En grupp på 5 pojkscouter står på en scen.
Tre unga pojkar spelar i en pjäs.
Två metallburar, den ena innehållande två kaniner, den andra innehållande kartonger.
Blå mjölk lådor sitter på en brygga vid en båt.
Två personer står på stranden en molnig dag poserar för kameran.
En man med glasögon som skriver på sin bärbara dator
Leverantörer sitter på en gatumarknad med burkar av varor som är röda och gröna.
En man i sjukhussäng med syrerör i näsan.
Två män, och en flicka bär flytvästar och simmar i vattnet.
En man är i en superbutik och handlar efter en Hawaiisk skjorta.
Två vuxna, två barn och två hundar sitter på en soffa.
En man i djup eftertanke medan kvinnan har mycket tålamod.
Fyra medelstora hundar brottas med varandra på ett gräsfält.
En flicka gömmer sig bakom en målad träkonstruktion inne i en byggnad.
En kvinna i vit klänning försöker ge en man i kostym kaninöron.
En ung pojke sitter i trappan med en bok.
En liten pojke tittar ut balkongen omgiven av växter, en leksak cykel, och plantera krukor.
En man cyklar med många olika föremål på sig.
En person som bär randig skjorta, blå jeans och blå gympaskor står på en sten i en bäck.
Två män på ett trafikljus som gör ansikten.
Två män som spelar bordtennis i ett rum med lägre belysning.
Männen sätter ihop metallramen.
En kvinna säljer grönsaker från en mobil gatuvagn.
En kvinna pratar på en mobiltelefon medan hon går längs en mans sida.
En person i gul skjorta pratar med en ung flicka.
Man med vit hjälm brinnande gummi av sin svarta och gröna motorcykel
En kvinna ser en brun hund springa iväg från ett hus tvärs över gräset.
En man som står framför en blå vägg och tittar ner medan han röker.
En man med paraply fotograferar under en mycket snöig dag.
Tre barn springer i ett fält runt cyklar
En ung man med glasögon, en svart skjorta och vit keps äter pizza och bröd.
En man kliver upp på ett steg från en trottoar.
En grupp på tre män och två kvinnor som sitter vid ett bord som har mat, dryck och ett spel på sig.
En liten flicka som täcker sina ögon i en gul skjorta, utomhus.
Två personer som kör motorcykel genom en mycket trång gata.
Parade utomhus med massor av ljus och färg.
En äldre kvinna som ser ut tar anteckningar i en föreläsningssal vid ett universitet, med yngre tittare studenter i bakgrunden.
En kvinna som sitter vid ett bord och tar en bild.
En man i svart rock ställer upp sin kamera för att ta bilder med.
Kvinnor i dräkter går över ett marmorgolv.
En man med vit hatt blir stampad av en brun häst.
Cowboy rider en häst medan två killar tittar från porten.
En man med ballonghatt håller upp färgade utskurna teckningar av två män.
Folk promenerar genom en inomhusmarknad.
En man står på trottoaren och håller en käpp i handen.
Folk fotograferar en byggnad.
En grupp människor är runt en hög med skräp.
En kvinna sår en indisk artefakt till en kommande festival.
En grupp människor i vita skyddsdräkter står framför svarta sopsäckar.
Två kvinnor tävlar i ett hinderevenemang.
Två unga mödrar besöker bordet vid matsalen och håller ett öga på sina barn.
En grupp människor tittar på en söt liten hund.
En kvinna i vit blus surar medan en man i svart skjorta tittar på.
En kille som jobbar i en fabrik.
En man på en tom trottoar nära en byggnad med en bakåt EC.
Ett barn gömmer sig under en möbel.
Folk står på en basketplan på en arena.
En ung flicka kysser sin mors läppar.
En svart man med röd mask bär en låda.
En ballerina klädd i gult är dans, på en scen.
En pojke i en röd poncho läser medan han lutar sig mot en stolpe.
Kvinna i svart promenader med barn förbi en väggmålning av ett torrt landskap.
En man med ett genomborrat ögonbryn tittar på en bärbar skärm, medan en katt är i bakgrunden.
Två rumskamrater försöker fixa diskhon i köket.
En dam i en röd mössa som serverar mat till samhället.
Två män i ett rum som pratar med varandra.
En man som ger sig i väg med händerna i ett rum fullt av datorer.
Man hjälper kvinnor med laptop i klassrummet.
Ett barn är ute och flyger med många ballonger i händerna.
En asiatisk man som står bredvid en dörr pekar på något.
En ung man står framför en grupp med några papper.
Man håller en bok och tittar bort från boken.
Unga kvinnor med päls och hatt går ut ur baren.
Någon lyfter en annan person på en karusell.
Två män spelar gitarr på scenen med två kvinnliga bakgrundssångare.
En man som förbereder en vit volkswagen att bogseras av en AAA-certifierad bogserbil.
En man i svart skjorta och en man i hatt uppträder på en konsert.
En kvinna som skär och säljer fisk.
En grupp unga vuxna som står inne i närheten av en ölutställning i Pabst Blue Ribbon.
En äldre gitarrist spelar gitarr på scenen.
En man och en ung pojke befinner sig i en flod nära en sandig strand.
Man med mörkblå förkläde tar en order
2 män med neutrala kläder har en konversation över en måltid.
En man som läser en tidning i en tvättomat.
Ett rum med asiatiska studenter arbetar i grupper vid skrivbord i ett klassrum.
En man med grå jacka och blå jeans talar in i en mikrofon medan han möter en publik.
En kvinna i röd utstyrsel joggar bredvid flera gatuskyltar.
Manlig gitarrist på scen i svart skjorta.
En man med mörk skjorta sitter bredvid en vit hatt och sover.
En person i en röd tröja seglar båt.
En ung kvinna med rött hår, klädd i lila håller i ett kuvert när hon går på en trottoar.
Flera människor som bär korgar på ryggen står bredvid varandra.
Unga vita människor sida i ett något mörkt rum.
En man i skinnjacka och cowboyhatt håller ut handen på gatan.
Ungt barn i en vit jacka som står framför en cykel.
Handske man som håller en rovfågel.
En man i lila kläder mjölkar renar med en skog i bakgrunden.
Killen tar en paus från att bära väskor upp trappor och njuter av en cup-o-noodles.
Två män, en bär gul skjorta och den andra en blå skjorta, spelar frisbee på ett plan.
Tre personer spelar frisbee i en park.
En kvinna som sitter i en solbränd stol bredvid en hund medan hon ler mot kameran.
Polisen griper någon på en livlig gata.
En ung man med LA på mössan målar en sköldpadda på en grön bakgrund.
En kvinna ställer sig i en sparkande position.
En man i vit och grå skjorta ser ut som en skjortlös man med mustasch rensar fisk på ett blekgrönt bord.
En patriot klär sig och sin häst med den amerikanska flaggans färger för en flashig uppvisning.
En brun hund hängande på en vit plyschleksak.
En kvinna cyklar på stranden.
En ung kvinna i en trenchcoat bär en plastpåse nerför trottoaren.
En vuxen och ett barn spelar monopol, barnet täcker sitt ansikte med handen.
Några människor går på stranden, skjutna från hög höjd
Människan sitter på toppen av balkongen och tittar på den vackra staden.
En kvinna i rosa bikini och en man i svarta badbyxor hoppar i vattnet på stranden.
En grön byggnad med två personer på framsidan.
En människa rider en häst nerför en grusstig.
Sandy beach, folk som går, ligger, sitter, en drake flyger.
En kock i svart skjorta och rutiga bandanna lagar mat på en industrispis.
En grupp på 4 personer gör olika aktiviteter från att spela gitarr till att använda en dator.
En cowboy på en knocking bronco i processen att kastas av ryggen.
Män i rinken med en man på utom kontroll häst.
En vattenskidåkare är luftburen ovanför vattnet nära en bakgrund av höga palmer.
En person som bär kappa och paraply är på väg hemifrån.
Mörke mannen använder en skruvmejsel för att bryta sig in i ett fönster i en gränd.
Två orientaliska personer sitter ett bord på en restaurang.
Tan färgade hund hoppar över en gren i skogen.
Två kvinnor äter middag tillsammans på en restaurang.
En man och en kvinna sitter nära varandra på en grön bänk.
En ung man som röker i en park.
En man lutar sig mot räcket på tredje våningen i en terminal.
En kvinna i gul skjorta på en tågstation.
Här är en bild på en tjej som bär en skjorta halvvägs upp och står bakom en kvinna som tittar ner.
Ett litet barn som får smak av dessertmix.
Ett litet barn i en rosa skjorta står vid en disk och blandar något i en skål.
En kvinna håller i en mikrofon när hon sjunger.
En afroamerikansk man, klädd i grön hatt, sitter utanför bredvid en koffert.
Fyra personer går nerför en gata, med två hålla händer och en hålla en gitarr.
En kvinna i brun jacka som skrattar åt nåt en vän säger till henne.
Två män på curlingarenan.
En man i röd kragetröja talar entusiastiskt in i en mikrofon.
Ett par står framför en tegelvägg som håller inköpspåsar.
En man i rött tittar in i ståndet hos en säljare på en marknad.
En man med rött skägg med grön Miller-hatt.
En kvinna i en grön tank övredel som håller en väska öppnar munnen och ser upphetsad ut.
En person med ett rött paraply som går nerför en snöig gata.
En man tvättar håret, borstar tänderna och rakar sig samtidigt.
En man går ut en lastbil medan han bär på möbler.
Många människor samlas för att titta på en ny uppfinning.
Kvinnan i blå byxor går förbi tegelväggen med graffiti.
En kvinna i svart beret och leopardtights sitter på en bänk.
Ungar väntar på paraden på gatan.
En kvinna i vit uniform sorterar nötter bakom en glasdisk.
En kvinna bär rosa tröja skära ost med kniv.
Fyra poliser står på en gata och en clown går framför dem.
Två damer klädda upp sig och festade på gatan.
Om utrustningen fungerar som den ska kan jag plocka upp varenda fläck.
En man på stolen annonserar eller delar med sig av information.
En man med randig svart och vit skjorta och hjälm rengör trägolvet medan en annan hjälper honom på bakgrunden.
En man väntar på att ta sig över korsningen.
Två äldre personer står på en trottoar med en hund i koppel.
Man sitter i en stol på ett utomhuscafé och röker en cigarett.
En snowboardåkare, klädd i en blå jacka och gröna byxor, snowboards nerför en kulle.
En man reflekterar under en stund vid en social sammankomst.
En brun hund simmar i det skumma vattnet.
En äldre man tar ett foto med en telefon.
Ett par klädda i vinterrockar beundrar inramade bilder på en vit vägg.
Religiösa män i bourgognekläder går nerför gatan.
En kvinna med cykel tittar på en staty, statyn är en display för en asiatisk restaurang.
En man skyfflar snö på trottoaren.
Två män pratar med en som tittar bort på avstånd.
En polis rider på en motorcykel på en stadsgata.
Flera människor sitter i en matsal med blått ljus ovanför dem.
En gymnast är balanserad upp och ner på en bar.
Runners, några i kostym, på en St Paddy's dag Marathon springa på gatorna som folk tittar på.
En kvinna håller i en bar medan hon tränar gymnastik.
En flicka i lila läder kramas av en tjej i blå och lila kläder.
En man går nerför en gata med cyklar bakom sig.
Två personer står ansikte mot ansikte på en bro nära en storstad.
Två män pratar som sett från ett skott.
En kvinna kramar en annan kvinna bakifrån.
Två personer har ett intimt samtal vid vägkanten.
En brunett i en skjortskjorta och knähöga strumpor, med gröna pärlor lindade runt handlederna.
Damen gräver genom sopcontainrar under en snöig dag.
En kvinna bär en morgonrock och bikini med klackar när hon står på scenen bredvid en blomkruka.
En kvinna går nerför en kall gata.
Här är hyreshusen och en försäljare som säljer glass utanför dem.
Kvinnor i rosa skjorta som säljer munkar i en park.
En man sitter medan han läser tidningen Times Sport.
Två personer går mot en person med tre miniatyrhästar.
En skulptur fungerar på en av hans verk.
En man promenerar längs en palmträdspromenad.
Två personer i kostym en grön en lila båda med vit ansiktsfärg.
Två ryska kvinnor pratar medan en tredje går förbi i förgrunden.
Två barn kramas medan de svingar ovanför en naturskön utsikt.
En kille i orange skjorta, orange skor och brun hatt på en luftburen skateboard.
Ett flygplan högt uppe i skyn med en man på marken.
Två personer gatustädning för hand och med maskin.
En man i grå rock går på en fallen trädstam i en skog.
En man sover på en röd bänk
Två personer organiserar en stor mängd mat utanför längs en livlig gata.
En person går förbi en gammal byggnad.
En vit hund håller en käpp i munnen medan den springer genom snön.
2 simmare i mitten av flyget gör ett dyk i en pool
En kvinna i en blå vinterjacka knuffar en kundvagn genom snön.
En kvinna delar ut flygblad till folk som går förbi.
En pojke som bär en röd "Jag älskar NY"-skjorta vinkar till någon till höger.
Folk går framför den utsmyckade tegelbyggnaden.
En man och en kvinna, båda i hattar, står på trottoaren i en upptagen stad.
En hemlös man med tjock jacka tittar på sin mat.
En kvinna i solglasögon och en hatt står på gatan med ett specialerbjudande smörgås ombord på henne.
En kvinna med glasögon som sitter nära toppen av en kulle och bredvid fordon för den terrängen.
En kvinna med svart jacka och röd halsduk och leggings går med en man medan en annan passerar och tittar tillbaka på dem.
En kvinna som står vid ett träd och tittar på sin telefon.
En liten pojke flinar i en folkmassa full av människor som poserar med slutna ögon i en sovande position.
En man i uniform står vid en ingång.
Två unga människor ler mot kameran medan de går sin hund.
En man hoppar när han snowboardar nerför ett berg.
En man och en kvinna, både i vita hattar, khakibyxor och mörka jackor korsar gatan.
En ung kvinna som går nerför de regniga gatorna i en röd parka.
En skylt finns i Times Square där man varnar för att Jesus snart kommer.
Pitcher är på väg att kasta bollen.
En person som vandrar vid foten av snötäckta berg.
En student som går på en trottoar nära ett campus.
En man sitter utanför vid ett träbord och läser en bok medan ankor äter i förgrunden.
En liten flicka i rosa kläder som håller gula stavar.
En liten pojke i en överdimensionerad mössa äter en isglass.
En grupp på fyra män går längs en strand, som en kvinna i en blå bikini ser på.
En man som bär en last av färska direkta lådor på bilen med hjul på stadens gator, när en kvinna går mot honom.
En man som korsar gatan under en kall vinterdag.
En ung flicka äter när hon sitter vid ett bord fullt av mat.
Man spelar in en video av en kvinna.
En kvinna i svart jacka som pratar i telefon i ett gathörn.
En äldre man läser en tidning på en trottoar.
Den här mannen bär en skjorta som säger "coolaste pappan i världen".
Vuxna som spelar fotboll utan uniform.
En flicka som bär röda shorts och sandaler sitter ute på ett räcke och flinar.
En kvinna som sitter i en stol och tittar in i en spegel.
En mörkhårig kvinna som får en vit klänning av en rödhårig kvinna.
En grupp unga vuxna som spelar Twister.
En kvinna med huvudband äter och en man ser på när hon äter.
En kvinna lägger nya matvaror på bordet.
Tre män sitter under ett blått tält på stolar.
En grupp människor står tillsammans och poserar för en bild.
Flera personer sitter på en bänk i ett offentligt rum.
En man sätter sig bredvid en rostig vägg.
Svart man sitter i förgrunden medan en mörkhyad kvinna i gul klänning går i bakgrunden med något i handen nära ansiktet.
En man i en smal allierad arbetar bredvid en affär medan en katt tittar på.
Flera män i rockar och jackor på en stad gata.
En man i en vit huva som håller en katt.
Folk passerar en hemlös person med en filt och röd huva på en isig gata.
En man som ivrigt trycker på i gräsklipparen på baksidan av ett hus.
En kvinna går med en barnvagn framför en byggnad.
Två äldre män som spelar fotboll med fyra barn som försöker göra mål.
Två män dricker öl framför ett stängsel.
En grupp människor sitter i gräsmattan stolar.
En gata är nästan öde med gul skylt öppnas upp bredvid en vit linje.
Folk står på en tågplattform under marken.
En kvinna läser uppmärksamt en tidning på tunnelbanan.
Bild av en asiatisk stad med människor som går längs trottoaren.
Två uppsatta poliser tar sig nerför gatan.
En cyklist närmar sig undersidan av en bro mellan byggnader.
En dam som bär en mörk dräkt och bär en vit väska går längs en gata.
Han går med en brun rock.
En man på en cykel med orange och svart tröja bär ett långt gäng pinnar.
En man med röd slips och kostym pratar med folk.
En ung flicka med en blå jacka kliver in i en pöl.
En man sitter och använder sin mobiltelefon.
En ung man i shorts som står under en trästruktur i grunt vatten.
Folk går längs en livlig stadsgata.
En kvinna som bär huvudduk går nerför gatan mot en infartsdörr.
Två fotbollslag tävlar på en fotbollsplan.
Kompakta bilar linjerar gatorna och en serie tält sätts upp längs en trottoar.
En kvinna går över trottoaren med 3 små flickor som håller varandra i handen.
En man och en kvinna undersöker noga en fiskespö tillsammans med en stor vattenförekomst.
En kvinna i svart klänning korsar gatan.
Ett klassrum fullt av barn som sitter vid blå skrivbord.
Folk står utanför nära en betongvägg och ett fönster.
En man i vit skjorta och blå jeans sitter vid vägen lifting, bakgrundsbildad av ett fält av blommor och ett stort grönt träd.
En kvinna i grönt hackar handen på en man i kostym.
En stor grupp människor står bakom ett podi på trappan till en kongressbyggnad.
Nancy Pelosi håller tal.
Två män och en kvinna sitter på en brun bänk med en brun hund.
En man vänder sig i luften inför en skara åskådare.
Fem personer, en man och fyra kvinnor, dras i en vagn av en mula en solig dag.
En stadsgata med en metallbänk upptagen av en kvinna i svart.
En skallig man kliver ur en liten blå bil.
En del människor går, sitter eller cyklar.
En liten flicka med en vit skjorta som spelar fiol.
Barn i ett grönt klassrum höjer sina händer.
En grupp svarta barn sitter bakom röda skrivbord i ett klassrum.
En skåpbil med flaggor reklam flyter, boogie styrelser, paraplyer, stolar och surfingbrädor.
Folk går på en livlig gata på vintern.
Två åsnor som drar i en kärra och bär gröna buskar, och de bär också människor på den.
Tre små barn i vita skjortor leker med en sten.
Ett barn som kör sin Power Wheels bil längs gatan, följt av sin pappa.
En äldre kvinna klädd i jacka, handskar och solglasögon knuffar en korg på en livlig stadsgata.
Två äldre kvinnor pratar med varandra.
Två män med hatt håller i sina cyklar.
Byggandet sker på en stor katedral.
Människan spelar piano utanför, med 3 observatörer, nära lyktstolpen, palmer och stora byggnad.
En polisman en New York-kyrka.
Tre personer går nerför gatan i ett asiatiskt samhälle.
Unga män spelar rugby på stranden.
Flera vuxna och en hund sitter på några vita stentrappor nära en grund pool
En blond kvinna tittar ner medan andra sitter i bakgrunden.
En man i cowboyhatt sitter ner och läser en bok.
En man i en skinnbiker jacka går trottoaren bär en stor ryggsäck.
En pojke ligger på en gräsbevuxen sluttning och en flicka står bredvid honom och läser.
Två brunettkvinnor i snygga, sexiga klänningar poserar för en bild.
En blond kvinna klädd i svart håller en kamera och stirrar på något på marken.
En vit bil står parkerad bredvid ett träd som har röd bark.
En man med hatt som håller två frisbee utanför.
En man och en kvinna pratar i en park
En ung asiatisk kvinna tittar på skärmen på sin mobiltelefon i en vit rock.
Två killar gör karaterörelser på en matta.
En brunett kvinna som bär en svart skinnjacka håller en lila handväska på en trottoar.
En man med bruna byxor RollerBlading.
En man med lockigt hår och skägg som går i folkmassan.
Välkommen till vår vackra plats och njut.
En man i öknen sitter på en häst som har massor av dekorationer.
En stor brasa brinner i skymningen.
Två damer går nerför en gata med svarta underkläder och gröna kjolar med strumpeband.
En man med hjälm som klättrar i ett snöigt område.
En rödhårig hona och brunhårig hane som bär glasögon promenerar tillsammans.
En folkmassa samlas utanför en vacker byggnad med en fontän.
Tre små pojkar tittar på kameran medan en av dem spelar på en hemmagjord trumma.
Flera unga kvinnor går nära blommande körsbärsträd.
En grupp ungdomar som går med två samtal på mobiler.
Två grupper av pojkar spelar en sport tillsammans med en boll
En grupp människor som korsar en gata i regnet håller ett paraply.
Fem personer och en röd telefonkiosk.
Tre personer står vid en vägg bredvid en vit byggnad
Två personer sitter i parken en kall vinterdag.
En man i overall och en hatt spelar akustisk gitarr utanför.
En fågel som sitter på en telefonlinje.
Två kvinnor joggar längs trottoaren framför en bensinstation.
En flicka i svart skjorta sitter ensam på marken.
En kvinna som bär solbränna är på väg ut ur en liten röd bil.
Folk slappnar av på cementtrappor med gräs, medan andra går förbi.
3 vänner som hänger i parken på gräset.
En gatuartist i vit skjorta och blå jeans drar i en publik.
Barnet är trött på den vandring han tog med sina föräldrar.
En blond kvinna i högklackat går förbi kyrkogården.
En man i orange skjorta framför bild på en man som håller i ansiktet och kramar ihop kinderna.
En liten pojke bär snorkel i ett badkar.
En svart man som stirrar på trottoaren med skuggor.
Flera personer står under ett klocktorn med två klockansikten.
En man i grå jacka och svart stickad hatt som går framför en grå upprullad garagedörr.
En man verkar sträcka sig efter en kvinnas drink på ett kontor.
En kvinna i lila topp och jeans pratar med en kvinna i en roller derby.
En person med en gul jacka som bär 3 apelsiner i en plastpåse.
Hon matar en get med getmat.
En blond kvinna lyssnar på hörlurar utanför.
En man i en vit trenchcoat med en väska som försöker ringa ett samtal på en telefonautomat.
En person som spelar dragspel på en bro.
En grupp människor och barn går längs en gångväg.
En man i infödingskläder passerar en skoaffär.
En kvinna, som bär shorts och en tanktopp, försöker skala ett rockansikte med hjälp av klätterutrustning.
En flicka handdukshänger sig på ett däck på stranden.
Det finns en person som står ett berg som har några intressanta former.
En get tittar på två pojkar precis utanför sin penna.
Ett litet gossebarn i GAP-skjorta sitter på en blå traktor.
Kvinnor står i dörröppningen på natten bredvid tågspår
En kvinna i svart njuter av det svala och uppfriskande vattenfallet.
En fotbollsspelare bär en grå skjorta och svarta byxor kastar en fotboll.
En man tittar på en TV-skärm i en restaurang.
En övergiven "Cafe Express" skylt är nu täckt av graffiti.
En man i hatt går i en stad och tittar åt vänster.
Kvällspendlarna går förbi bussar som kantar en stadsgata.
En man sitter i en båt med två andra män som paddlar vattnet.
En man och en kvinna stirrar på ingången till några katakomber.
Två män bär vita skjortor med hjälm när de cyklar.
En man med smutsiga kläder sover på trottoaren.
Ett gäng barn i kanoter på en flod.
Fyra kvinnor är utanför en kinesisk affär.
Folk cyklar bredvid en blå och grön buss.
Mannen som låg på ett delvis byggt hus.
En kvinna i rutiga byxor står på en skidbacke, redo att gå ner.
En läkare tröstar en idrottsspelare skadad.
En man och två kvinnor som äter och dricker i ett kök.
Pojkar i uniform väntar utanför en byggnad.
En äldre kvinna i en kappa som går nerför gatan.
En gammal kvinna med en käpp som går bredvid en bil.
En man som tittar över balkongen i en modern byggnad.
Två flickor i gröna tröjor poserar utanför.
En grupp människor som går tvärs över gatan några bär stora svarta och röda flaggor.
Den åldriga kvinnan sitter medan hon bär sina rosa-linsade glasögon.
En grupp barn är ute klädda i blått i ett inhägnat område.
Folk stirrar på marknaden.
En pojke i en blå jacka pekar ut något för sin mor, också bär en jacka, när de går igenom en färgstark karneval scen.
Ett litet barn som ligger på ett trägolv.
En rad röda cyklar står parkerade på gatan.
Ett barn ställer sitt huvud genom ett hål i en målad vägg.
Två män fotograferar rosa blommor, en med en liten digitalkamera och en med en större lins.
En liten pittoresk stad som alla lyste upp under semestern.
Person i röd hatt som går på trottoaren en snöig dag.
En äldre man spelar saxofon.
Mannen med rakat huvud och skägg poserar på en expansiv strand med en orange sandhink på huvudet.
En byggnadsarbetare blåser skräp från trottoaren
En man, klädd i vitt, håller en burk medan han går på tegelsten.
En man i grön jacka spelar en fairground spel.
En kvinna i blå jacka går bredvid en affisch med två gröna figurer som ser ut som män.
Den svarta och bruna hunden springer genom snön.
De som letar efter män hänger vid vägkanten.
Mannen i brun kostym går mot kameran nära raden av bilar.
Instrumentbrädan i en bil med en brun hundleksak och en rosa docka.
En man i jacka sitter och snokar på en grön parkbänk.
En man och en ung blond pojke som använder interaktiva plastleksaker utanför.
En flicka sjunger medan hon hoppar i luften.
Ett par som var täckta av färg fångade uppmärksamheten hos dem som stod framför dem vid fruktstället.
En amerikansk postlåda täckt av graffiti.
Män i turbaner tittar på medan man greppar en kamel vid halsen.
Unge man jobbar hårt vid sjön.
En kvinna går i snön med en polka prick paraply.
Tre män går på en trottoar i en stad.
Tre arbetare går ut ur sin säkrade byggnad i slutet av dagen.
Kvinna med rosa skjorta sitter i stolen.
En kvinna med en svart väska som går ut på gatan medan en man i kostym går till vänster.
En man talar en presentation medan andra tittar på ett bildspel.
Killen i mörk kostym på podiet pekar mot powerpoint-skärmen.
En limousin som kör nerför en gata i ett graffiti-laten område.
En närbild av en kvinna som går medan hon bär en svart och blå tanktopp med solglasögon ovanpå huvudet.
En kvinna som står på trottoaren med händerna i fickorna.
En grupp människor passerar genom torget.
Flera vuxna går nerför en stenlagd gångväg i Europa.
En person som knuffar bagage och någon på mobilen i en stad.
En gammal kvinna på en kall dag, utanför en sportaffär någonstans i Brasilien.
En kvinna i solglasögon står bredvid en orange skylt som läser RoadWork Ahead.
En man i en stad går över gatan och kör en kärra.
Tre unga pojkar är klädda i hoodies vända på samma sätt.
En man som håller sig på gatan och tittar bort från en tiggare.
En man med ryggsäck går nerför trottoaren framför en röd tegelbyggnad.
En kvinna i en vit tanktopp går och håller något i sina händer.
Fyra personer, tre män och en kvinna, arbetar på sina datorer.
En polis med hög siktväst håller en stoppskylt.
En kvinna som bär svart bär en behållare med mat.
Ett äldre par läser en karta på en parkbänk.
En gammal man i rock och hatt sitter på en parkbänk.
De här kvinnorna tittar på när folk spelar tennis från en bänk.
En kiteboardåkare som bär hjälm och glasögon rider över ett snöigt landskap.
Två små barn tittar på färsk hummer i mataffären.
En man i rött går framför en vägg av fönster.
En kvinna som sitter i en tågvagn.
En cyklist som väntar på att trafiken ska passera så att han kan korsa gatan.
Ett litet barn som leker på ett dammigt torg.
En kvinna håller en frusen pop sickle och nycklar i sin högra hand.
Två kvinnor går runt i en stad.
En man i uniform sitter på en stol med ett gevär vid sin sida.
Gammal kvinna i vit skära färgglada hantverk som lakan.
En äldre kvinna med käpp går med ett tecken runt halsen.
En man målar en bild på trottoaren.
Äldre kvinna går nerför stadens trottoar i en gul jacka som håller en svart Zales väska.
En kvinna som sitter vid en soptunna.
En medelålders man läser tidningen och dricker Starbucks kaffe i parken.
En gammal man på ett tåg läser en tidning.
En man i svart jacka som sitter på en buss med hörlurar.
En gatuförsäljare med mörkt hår och glasögon, sitter på en fällbar stol.
Några personer går på avstånd från en liten stad.
En man knuffar en cykeldriven vagn nerför tegelgatan.
Tre manliga studenter arbetar i ett labb med en av dem tittar genom ett mikroskop.
En grupp vänner som går längs trottoaren.
Tre kvinnor tittar tillbaka på kameran som sitter i baksätet på en skåpbil när föraren kör längs vägen.
En rödhårig kvinna i svart rock framför ett tecken.
En äldre man i svart jacka och blå jeans sitter på en bänk medan han tittar på sin telefon.
En kvinna läser en tidskrift medan hon sitter vid ett bord.
En ung man på en fest skriker ut, hans knytnävar lyfts av känslor.
Två bruna hundars råa hus utanför.
En äldre man klipper håret på en kund i sin frisörbutik med blomsterväggar.
En man i röd jacka ler när han håller en cykel över huvudet.
En man i blå skjorta ligger på stenar i solen.
En kvinna talar in i en mikrofon vid en social sammankomst.
Många bilar på gatan, och en man på cykeln.
En äldre kvinna cyklar tvärs över gatan framför en stor grön byggnad.
En attraktiv ung dam ute i offentligheten glänser i sidled på något utanför kameran.
Flera män och kvinnor samlas på ett idrottsevenemang.
En vagn med paraply sitter mellan två män.
En man i röd jacka och hjälm cyklar.
En afroamerikansk manlig ungdom rider en grön cykel medan andra människor tittar på bilder på en bräda.
En bil får böter för en parkeringsintrång.
En indianfamilj står tillsammans, djupt i en vattensamling och ser upp.
Fyra musiker som spelar gitarr på en klubb.
En man med en gul hatt på lutar sig mot en vägg av något slag.
Flera personer går upp för en uppsättning utomhustrappor.
Ett barn i svart rock löper över en graffititäckt bro.
Två personer står i en blomsteraffär.
En man går 11 hundar samtidigt.
En trio med tjejer klädda för att gå på fest
En sittande kvinna skrattar bredvid en man i en blå jacka.
Barn som sitter på sten i öknen
En grupp pojkar som bär ärmlösa vita skjortor dricker ur en vit kopp.
En blond tjej och brunetttjej som går.
Tre män jobbar på ett tak, medan en man klättrar uppför stegen.
En ung pojke arbetar jorden på sin gård.
En man med svart hatt går med en klyfta.
Glad mamma vänder sin dotter runt och både leende öra till öra.
En hane och en hona i lätt färgade kläder dansar.
Medelålders man, med skinnjacka, står på en dimmig parkeringsplats.
Volontärer är på den här bilden med sin hund som letar efter en saknad flicka som senast spelade i skogen.
En skolös ung pojke sitter på toppen av en stenhög.
En äldre kvinna, en yngre kvinna, en ung pojke och en svart pälshund som går på en grusväg i en skog.
En kvinna och en pojke njuter av en promenad i skogen.
En kvinna och ett yngre barn går i skogen.
En kvinna som går förbi en minibuss och husbil i skogen.
Barn leker på en lekplats uppsättning med varandra.
En man klädd i inbördeskrigskläder har en musköt.
En konstnär som bär en röd gingham scarf arbetar på en målning av ett torn.
En flicka i rosa hatt sitter på marken.
En kvinna går förbi en garagedörr som säger "ingen parkering när som helst".
En pojke som skateboardar nerför en brant lutning.
Mannen i röd skjorta och blå jeans justerar sin fluga.
En man som går i en vit morgonrock.
Två stora män är klädda i svarta t-shirts, khaki bottnar, stövlar och smycken med hårdvara.
En man spelar musik med svärd och båge.
Mannen i den röda skjortan låtsas spela fiol med ett paraply.
En kvinna med en stor väska och stövlar som går i en marmorliknande hall.
Två hundar med skjortor leker i det gröna gräset.
Två cyklister tävlar nerför en gata.
En man och en kvinna sitter på en bänk.
Fyra personer går genom en stad.
Folk springer i någon sorts maraton medan de passerar blå skyltar.
En kvinna i grå klänning går.
Tre tjejer går nerför gatan medan den i mitten studsar en svart basketboll.
En man i orange rock sitter på en motorcykels passagerarsäte.
Fyra personer går ner från eltrappan, klädda i väldigt varma kläder.
En grupp människor äter lunch i ett fullsatt café.
Ett barn i en vit huva springer mot en flock vita fåglar.
Ett par som håller varandra i handen går nerför en gata.
En kvinna i svart med ett rött paraply går mot en katedral på en asfalterad gata.
En kvinna knuffar en pojke i en vagn nära en trottoar.
En man i blå jeans målar en väggmålning på en ljusblå bakgrund.
Folk samlades vid ett utomhusevenemang.
En kvinna som sitter vid ett bord och tittar noga på sin Apple laptop-skärm.
Par av kvinnor som håller parasoller går nerför en gata i vått väder.
Person i en blå anorak som läser en stor skylt stående på en tågplattform.
En Santa Cruz brandkår motor utanför en Gap butik.
En ledsen liten pojke som sitter vid ett bord med en blå duk och äter chokladglass.
En grupp bilar, bussar och cyklar täpper igen en gata.
Fyra personer med skotrar framför en mycket stor metallport.
En kvinna som håller i ett gult paraply i regnet.
Här är en tjej i stövlar som går med ryggsäcken under ett paraply i regnet.
En skjortlös, tatuerad man med hat bär en skateboard.
Restaurangpersonalen håller på att sätta upp matsalen för en måltid.
En äldre gentlemän i rött går förbi en person som bär allt blått.
Två barn, en i röd jacka och en i blå jacka, sitter i en däcksvinge.
En läkare med sina assistenter arbetar under ett tält.
En grupp läkare samlas runt en patient i ett operationsrum.
En afroamerikansk kvinna som bar gul frukt på huvudet och gick bort från en byggnad.
Två kvinnor, en i blå skjorta och en i grön skjorta, går över en livlig gata med kastruller på huvudet.
En blond kvinna bär en jacka med ett öga på den.
Fotgängare bombarderar en stad gata täckt av konsumism, inklusive skyltar för Burger King, McDonalds, Subway, och Heineken.
En hund hoppar och fångar en blå boll i munnen.
Kvinnan i den lila bikinin och rosa övredelen bär en hjälm.
En fullsatt stadsgata med många fotgängare.
En kvinna i brun tröja och jeans tar en bild av en kille med skägg medan en annan kvinna sms:ar på sin telefon i närheten.
En person sitter på en stol medan han lyssnar på musik.
En skräckslagen fotograf i kostym tar bilder av en grupp små barn som sitter på marken.
Hunden springer med en lila leksak i det snöiga fältet.
En man i en T-shirt spelar schack.
En man bär en sopsäck tillsammans med sin käpp.
Två personer på en cykel bär stora hjälmar med personen i ryggen klädd i lila stående på fotstöd på baksidan av cykeln.
En man i gul skyddsjacka och blå jeans sitter på mobilen.
En kvinna som håller en gul väska framför en "Välkommen till Aberdeen"-skylt.
En äldre hane jobbar på en snöbil.
En kvinna med en kamera som många bakom henne går över vattnet på en gångväg.
Barnens skidklass är inställd på att lyssna på instruktören.
En kvinna går nerför en gata med ett paraply.
En kvinna som målar med en rulle.
En man och en kvinna sitter utanför - Kvinnan bär päls och mannen ser professionell ut med slips.
En man som kör motorcykel i sidled i Japan.
Ett litet barn som bär en rosa jacka med huva och orange byxor springer.
En grupp hiply klädda unga vuxna slappnar av tillsammans.
En pojke som leker i vågorna, med en mås i förgrunden.
En man i svart som går nerför trottoaren och tittar på sin I-Pod.
En man läser en tidning sittandes i ett tåg.
Två män går längs gatan och går åt motsatt håll.
En kvinna poserar med ett barn i bakgrunden som leker med bubblor.
En man som står i ett stort rum vid ett fönster.
Kvinnan i vit hatt och blå cape står nära shoppingvagnen på en livlig gata.
En ung kvinna med beige byxor går en hund.
Bilar kör under en bro medan folk går upp.
Ett ungt indiskt barn håller en docka längs ett staket.
En man i grön tröja pratar i telefon och håller en flicka i knät.
En kvinna i en ytterrock använder sin telefon när hon står utanför en byggnad.
Unga par tittar på en butiksutställning under ett paraply i regnet.
Följer du med mig på en kopp kaffe?
Tre personer i en linje som korsar en gata framför en delikatess.
Den här personen gör glasstrutar.
Flera människor går medan de bär rockar, medan man cyklar.
Det finns 6 vänner som går nerför gatan.
Två personer i lila kyss bredvid ett provisoriska tält och camping.
En grupp människor samtalar med varandra.
2 man och en hund går nerför en väg bredvid fält
En byggnadsarbetare flyttar en apparat utmed en räls framför en byggarbetsplats.
En person äter en tallrik pasta med en svart och brun hund i knät.
En man som kör en scooter längs en kullerstensväg.
En man och pojke sitter korsbenta på marken och inspekterar grillen.
En man går förbi en dieselpåfyllningsstation.
En kvinna i en grön blus står på vägen och tittar på mörka moln som samlas på avstånd.
En man på gatan som ritar bilder av människor.
En ung svart kvinna har en skylt som erbjuder fria kramar bland en skara människor.
En pojke i röd skjorta och jeans försökte röra motorsågen.
En man hoppar med sin cykel på en parkeringsplats bredvid en fyrvåningsbyggnad.
Två kvinnor pratar med en okänd person på en trottoar.
En man med röd plastnäsa och randig tröja som håller i en glaskula.
Två kvinnor håller rumpan av en naken man
En man i glasögon bär en mörk rock.
En man i röd skjorta som kissar utanför vid ett träd.
Människor som sitter på en lägre nivå av en gångväg, medan en annan person går ovanför dem bland träden.
En gammal man med glasögon håller i en pinne.
En grupp människor som sitter vid ett bord och äter.
En svart kvinna med flanelljacka och papperspåse går nerför gatan.
En kvinna som läser en bok på en bänk i en park.
En äldre man i blå skjorta lagar mat.
En man i grön jacka med glasögon bär en massa blommor.
En parkeringsplats med en cyklist som rider genom den.
En man står mitt på en väg och pratar på sin mobil.
En kvinna håller gröna och guld pompoms.
En förvirrad man står och stirrar ut i fjärran framför några biljettinsamlingsmaskiner.
En man och hans tjej går över gatan.
En person med blå hjälm på med svarta stövlar, som rider på en häst.
En man sitter på ett kontor och tittar på en datorskärm.
En kvinna i svart jacka och en svartvit randig kjol tittar på en kvinna som pratar med en liten pojke som sitter på betongtrappor.
Shoppers går på en upptagen stad gata.
En kvinna i grå rock, med brunt hår, drar en korgliknande vagn.
En person rider havets vågor.
En man väntar vid en busshållplats med en rosa fyr och en grön båt i bakgrunden.
En hund sprutas med vatten i ansiktet utomhus.
En mor och hennes två barn framför en gammal, sliten byggnad.
En hund går ensam på ett fält.
En ung man på en segelskida som bär en torr kostym mitt i en vattenförekomst
Grupp av hundar som går och sniffar på grus.
En yngre kvinna som sitter nära en vattensamling med en hund.
En ung man i solglasögon tar en paus från sitt jobb.
En kvinna i blå topp och pennkjol går förbi en flintskallig man i en spetsig kostym.
En man i blå kostym går nerför gatan.
En man i en diamanttryckt tröja och jeans står mitt på en trottoar och lyssnar på öronhandtag.
En kvinna med en gul väska springer över en livlig gata.
En man klädd i svart står vid ett gathörn nära ett korsande ljus.
En ung kvinna i blå Hollisterskjorta och blå jeans.
Tre män med hattar sitter och dricker vid ett bord.
En kvinna som är upptagen med att multitasking på telefon och dator.
En vit cykel är bunden till en gatuskylt.
En flicka är koncentrerad läsning på sin eReader.
En man sitter på en bänk med sin cykel utanför staden.
En kvinna som pratar på en mobiltelefon och håller i ett paraply.
En pojke i blå skjorta plockar upp något från marken medan en publik samlas.
En man sitter och håller fram en kopp.
En kvinna sitter på vägen bredvid sin cykel.
En kvinna i svart och en jeep i blått.
Fem barn leker i en översvämmad (eller avsiktligt vattnad) lekplats.
En blondhårig kvinna spelar dart i en bar.
En äldre kvinna som bär solglasögon tittar genom sin handväska på en fullsatt marknadsplats.
En kvinna går över en veranda med en yxa.
En grupp män i vitt, blått och svart marscherar ut med ett jättekors.
En spansk man som bär radband väntar på en taxi.
En kvinnlig barista som bär svart gör kaffe i ett kafé.
En ung pojke och mörkhårig man tar bilder i motsatta riktningar.
En hund springer genom ett fält med tungan hängande ut.
En långhårig kvinna lutar sig mot ett stenräcke och tittar ut över havet.
En liten pojke i en blå hjälm som leker med en gul leksaksbil.
En grupp människor går genom en tunnel.
Fyra personer är i en paviljong och får drinkar av två män.
Två personer går på en randig stig.
En person rider en fyrhjuling genom ett lerfält som har flera byggnader bakom sig.
En tjej kastar en softball till sin lagmedlem på basen.
En ung man med lila hatt skrattar med tuggummi i munnen.
En man och en kvinna står vid skylten.
En medelålders man får huvudet helt rakat av en annan medelålders man med hår.
De är här för att se till att ingen korsar barriärerna.
En man klädd i svarta samtal med en dam klädd i en ljusblå klänning och en vit huvudduk.
En man som kör en kärra dras av en åsna.
Pojke, ungefär 10 år gammal, som ramlar ner i en orörd pool på en varm sommardag.
Två män står och ro en tunn båt i havet.
Två personer går runt på en livlig gata.
En man som spelar dragspel rider tunnelbanan i New York.
En man som går in i en byggnad när en annan man sitter på en gata en kall dag.
Folk förbereder sig för ett modellplansmöte.
En dutchfamilj samlas runt ett påskägg som består av blommor.
En man serverar mat vid ett matstånd.
Ett kvinnligt barn som bär en rosa skjorta leker på en lekplats.
I en skog diskuterar en man och en kvinna något.
Män i soldatuniform skjuter vapen i luften.
En liten hund som tuggar på en svart rem.
En kvinna i blå kläder ler när folk i bakgrunden går förbi.
En kvinna klädd som sjöjungfru Ariel bredvid en telefonkiosk.
Två kvinnor i kostym, den ena klädd som sjöjungfru, den andra som älva, delar ut broschyrer.
En liten flicka som sitter på en bänk med en boll under.
En man i vit skjorta går hand i hand med en kvinna som också bär vitt.
En clown i en röd spetsig hatt som skapar ballongkonst.
En kvinna i en rosa tröja som sitter bredvid en man i en vit vindjacka framför en mobil matbil.
Man med sjal ber vid en stor sjö och liten båt.
En kvinna klädd som en sjöjungfru i en lila snäckbh ser till vänster.
En kvinna sover bakom disken i en affär.
Tre män sitter bredvid varandra och mannen i mitten läser en bok.
Sex personer på en klippa tar en bild av deras vatten.
En man i en rosa och vit randig skjorta som håller en hästs tyglar.
En kvinna som går, bär en skogasmväska.
En man arbetar med eld och tjära för att reparera ett tak.
Två personer med baseballtröjor som hoppar i luften.
En ung man cyklar på en yta täckt av graffiti.
En jonglör som sitter för sig själv och jonglerar med bowlingpinnar.
En pojke sitter i en barnvagn med en blå hatt och röda vantar på.
Folk lutar sig mot att bevaka stan.
En man i rutig skjorta sjunger och spelar gitarr.
En kvinna spelar gitarr.
En ung pojke i svarta byxor och en blå skjorta har just sparkat en fotboll.
En kvinna tittar in i fönstret på ett franskt bageri.
En äldre kvinna med brunt hår går sin cykel genom en grind till en trädgård.
Förbudet i den svarta hatten är att leka charader med sin vän.
En man som bär svart och svart hatt häller en dryck i en kopp.
Ett par som ser ut som om de är förälskade.
Det finns 5 män i en liten motorbåt, bakom dem finns en tropisk djungel.
En man och kvinna rider i en mulåsna dragen vagn som föraren pekar ut landmärken.
Mannen i mitten lyfter armarna när han och de två kvinnorna möter podiet.
En man och två kvinnor sitter på en bänk.
Ett barn står tillsammans med en äldre kvinna vid tunnelbanestationen 96th Street.
Folk glider ner för en jättegul och röd rutschkana.
En kvinna med hörlurar i öronen går nerför gatan medan en man som pratar på sin mobil går bakom henne.
De tre flickorna uppträder någon form av dans.
En tjej i en röd rutig skjorta med blå jeans som gör en knytnäve.
En flicka hoppar på gatan på natten medan en annan flicka tittar.
En person som bär en blå och gul snödräkt, en blå hjälm och snöglasögon rör sig nerför en snötäckt lutning.
Två pojkar står framför varuautomaterna.
En rynkande äldre person går och bär en plastpåse
En kvinna och en man som sitter på en soffa i en affär.
En rödhårig kvinna sitter på en soffa med korsade ben.
En grupp afrikanska män lastar en lastbil full av färsk fisk.
En man i vit hatt står på gatan och håller färggrant papper.
Två män spelar instrument på trottoaren.
En långhårig kvinna klädd i keps, jeans och gul skjorta verkar leda en osynlig hund med en förlängningsbar koppel.
Ett par asiatiska människor äter glasstrutar.
En man i grå jacka spelar piano på trottoaren.
Två tonåringar stirrar över ett bord.
Ett ungt par går längs en bäck en varm dag.
En man i grå t-shirt och jeans hoppar i ett vardagsrum.
En man med en klipphök håller flera trämöbler i ett plastbad i gathörnet.
En tjej i bikini tar en bild av några personer.
De som står på Washington Wells-plattformen och väntar på ett tåg.
En idrottsman bär neongröna och orange snowboards över en liten blå bil.
Två hanar går medan en hona håller i ett paraply med vita prickar.
Flera byggnadsarbetare som står på en ställning
En nyfödd pojke ligger i en inkubator med många rör.
En ung person gör ett trick på en cykel.
Ett par poserar med sina snowboards mitt i ett snöigt virke.
Blå halvbil och två herrar som står framför den.
En kvinna med genomborrad näsa är under ett blått paraply.
En man i svart rock går.
En gul bil kör genom gatan med tre fotgängare på en trottoar.
En man som bär många påsar burkar kommer förmodligen att sälja dem för skrot.
En kvinnas hand och arm med blå naglar och en tatuering som inte är ångerfull.
Ung flicka med målat ansikte och flätor sitter på en bänk vid vattenbrynet.
En herre i en keps skriver böcker åt ett par kvinnor.
Den här tjejen är klädd i en röd snödräkt och klättrar i ett träd.
Efter att ha fallit ner i snön tar en ung kvinna ett foto av sina vänner på avstånd.
En man som står bredvid gatan med gitarr på ryggen.
En mycket lång kvinna i en mycket kort orange klänning promenerar nerför en tom trottoar.
En pojke med väldigt ljusa gröna luddiga byxor.
En blond kvinna skrattar åt kvinnorna bredvid henne med en vit fransjacka.
Två honor som springer runt på ett spår, i idrottskläder.
En tatuerad man som städar rännstenen med en spade.
En person går framför helarens affär.
En kvinna klädd i svart topp och grön kjol dans, som en man i bakgrunden ser på.
En liten flicka sitter på huk bredvid en vattensamling medan hon petar en käpp i den.
Två personer i rockar som går bredvid ett staket.
En man som väntar på bussen i ett krigshärjat land.
En person som bär en brun huvtröja och jeans med ryggsäck går nerför gatan.
En kvinna i tunnelbanan tittar ut genom fönstret.
En man och en kvinna som ligger på röda metallbänkar framför en stads skyline en solig dag.
En ung kvinna som bär huvudduk går nerför gatan och bär sin handväska.
En kund i svart jacka tittar på fina ostar.
En fotbollsspelare sparkar bollen.
Folk sitter i läktarna på ett idrottsevenemang medan andra står ut på spelplanen.
Han gör sig redo att sparka bollen.
En man i hatt och rock pratar i telefonen bredvid en byggnad med ett tecken som är på ett främmande språk.
En man knuffar en docka med några lådor nerför en stadsgata.
En man går över en gata med sin son.
En man och en kvinna som omfamnar på trottoaren.
En kvinna i skinnjacka gäspar när hon går bredvid en ung pojke på trottoaren.
En biker, klädd i svart, går längs en väg till sin cykel.
Athlete i svarta shorts som springer nerför en trädkantad gata.
En man på en cykel rider förbi en man och hans son.
En gammal man sträcker sig efter sin frus hand när de går över gatan.
En kvinna och ett barn som korsar gatan.
En man i svart keps och jacka sitter på blå väska framför en byggnad.
En äldre kvinna som håller i sin handväska medan hon beundrar många ljus.
En kvinna i en röd tröja står bredvid lådor med ananas.
En äldre man i kostym som drar sitt bagage bakom sig.
En flicka i en blå halsduk och grön skjorta står bredvid en röd cykel.
Två killar spelar i ett band, en spelar gitarr och en spelar tangentbordet.
En smal skateboardåkare hoppar över en brandpost på sin skateboard.
Människor samlades kollektivt för att hedra ett ögonblick i tiden.
En stor grupp människor samlas framför en hög byggnad.
Ett barn i hatt och jacka tittar på blommor.
Man med kort hår i en blå jacka tar ett foto av en stor grupp människor som står framför en stor upplyst byggnad.
Ett nygift par står nära en bil.
Titta noga när jag visar konsten att glida en frisbee.
Tre killar uppträder i ett band på scenen.
En man utför stunts framför en publik på trottoaren.
En akrobatisk underhållargrupp demonstrerar för intresserade åskådare.
Flera män och kvinnor sitter runt i en hydda och väntar på att deras tur ska bli nästa.
En kille som visar sin cykel för ett barn.
En man i vit skjorta sitter framför en mikrofon och spelar gitarr.
En man i svart skjorta spelar gitarr.
Flera människor bär färgglada kläder och hattar presterar i ett öppet område.
En man i blå overall hänger på en stolpe ovanför en folkmassa.
Personen i en röd mössa tittar över vattnet medan han sitter på en träbänk.
Ett par tar med sig hundar på en promenad genom parken.
En man i urban gatuutrustning med en randig huvtröja tittar ner på något i sin hand, framför en tegel-och-glas butiksfront.
Det finns en bro över en vacker scen av byggnader och vatten.
En man går en orange hund framför en byggnad med ett rostat kedjestängsel.
En far med sin son på axlarna som går genom en park.
En äldre man säljer tidskrifter i en tidningskiosk i Asien.
En man sjunger i kyrkan.
En man går över en gata på en solig dag.
En skjortlös kille vände sig om och filmade något på stranden.
En kvinna i lila topp står i ett rum med en röd vägg.
En kvinna ritar en karikatyr av en ung pojke.
En man sitter på en parkbänk och tittar på vattnet.
Man i grå och blå rock blåser bubblor.
Kvinnan med brunt hår och vit rock står vid skylten "Shine Deli".
En snowboardåkare på en bergstopp i en klargrön jacka.
En man och kvinna tittar på en karta i Central Park.
En dam bär en gråtande pojke på trottoaren.
Tre barn ställde upp för att få mat vid ett bord.
En kvinna i en brun tröja justerar sina glasögon.
En valp utan svans hålls av sin krage av ägaren.
En målare sätter eftertryck på en bild.
Två unga pojkar som spelar lacrosse springa för lacrosse bollen.
En kvinna är på väg ner på rulltrappan.
En kvinna pekar nerför gatan till sin vän framför en ingång till en tunnelbanestation.
En far och son som leker med ett trätåg på en stadsmatta.
En man i röd uniform står utanför Broad St Station och pratar på en mobiltelefon.
Skäggig man med strumpor med sandaler sittande på en bänk.
En kvinna skjuter en skottkärra medan två andra tittar på i en park
En pojke kramar en mindre pojke bakifrån.
En äldre person mot en vägg på gatorna tittar ner med en kopp och fotograferar i handen.
Två små lacrossespelare lyssnar som de instrueras.
En man med gitarr framför en grupp tjejer med hattar.
Tjejer i kostymer som pratar med säkerhetsvakter.
Fyra flickor i röda uniformer bestående av röda tröjor och röda kjolar går nerför gatan.
Män och kvinnor i färgglada kostymer dansar.
Två kvinnor som bär halsdukar på huvudet joggar på ett strandbad.
En kvinna säljer handgjorda hattar.
En man i grå skjorta som spelar röd gitarr.
En man spelar gitarr medan en annan man fotograferar.
En stor hund hoppar över ett fallet träd i skogen.
En grupp män som spelar och sjunger musik medan en publik tittar.
Två män på cyklar passerar en rad byggnader som specialiserat sig på medicinska tjänster.
Ett gult tåg är på spåret.
Två kvinnor står utanför och tittar på något med roliga uttryck i ansiktet medan de andra människorna omkring dem inte verkar märka det.
Någon med en orange jacka som går med en cykel pekar mot en byggnad.
Tre barn ler framför en annons för en kamera.
En man ger en liten flicka en puss.
Denna bild är tagen utanför och har en ung flicka tittar med ren glädje som hennes pappa visslar till henne.
En elev får hjälp med läxorna.
En grupp barn som leker i en vattenfontän i sina badkläder.
Vägarbetaren bevakar en inkommande cementbil.
En surfare går längs stranden när han ser ut över vattnet.
En man i alla blå kläder som paddlar kanot ensam.
Fiskare kastade nät från utgrävda kanoter i vattnet.
Tre pojkar håller uppblåsta cykeldäckringar på en dammig stig.
En man i hatt står bakom en gatuuppvisning av solglasögon.
Två personer och ett barn som går genom en flod.
Pitcher i ett basebollspel med en vit 34 uniform som gör sig redo att kasta bollen.
Fyra kvinnor och en man spelar kinesiska pjäser i någons hem.
Bara ett fåtal människor njuter av dagen på stranden nära den gula bulldozer.
En liten flicka som ler lyfts upp av en vuxen.
En kvinna i röd jacka dricker på motorhuven på en bil.
En man med en kamera som stirrar på en staty.
Folk svingar på en gunga i en park utanför flera hyreshus.
En ung man som åker skateboard över en ramp bakom ett kedjelänkstängsel med två vänner.
Två kvinnor går på gatan hand i hand på natten.
Det finns en man i glasögon och en labbrock.
En man och en kvinna sitter på en picknickfilt på ett fält ett grönt gräs.
En blond man i brun läderjacka lyssnar på musik.
En baseballspelare springer till en bas, medan hans lagkamrat glider till en bas i bakgrunden.
En basebollfångare är redo att kasta medan hans lag tittar på.
En flicka stänker vatten i en pickup som kör förbi.
Tre kvinnor står utanför en byggnad och pratar med en man.
En kvinna poserar framför ett kuperat landskap medan hon håller i ett träd.
En man sitter på en bänk med en vit hund i närheten.
En rad börjar bildas på The Cheap Tab Shop.
Ett par honor pratar med varandra medan en snärtar sin cigarett.
En man i rutig röd skjorta kastar ut sin fiskelina i vattnet.
Barn bygger sandslott på stranden.
En afrikan som kikade ut ur ett tunnelbanetåg i New York vid Wall Street-stationen.
En man och en kvinna står vid en parkeringsplats och pratar på mobiler.
En kinesisk kvinna med hål i jeansen pratar på en mobiltelefon.
En affärsman som går på en gata.
En blond kvinna står ensam i en gränd.
En ung kvinna i jeans går nerför en gata.
En vit man i telefon och en svart man som sitter i vita stolar.
En man i orange skjorta som tittar på sin mobil.
En kvinna lämnar en tunnelbanestation medan hon lyssnar på musik.
Två män klättrar uppför en trappa.
Två män med hårda hattar är på en arbetsplats.
En förlorad hund som försöker hitta mat på en pizzarestaurang.
En stadsgata med ett hål i mitten.
En man i röd tröja väntar på ett gatukök.
En elektriker observeras från ett fågelperspektiv som arbetar på en transformatorlåda.
Alla dessa människor väntar på att gå över gatan.
En tjej som dansar mitt i en grupp människor i parken.
Tre kvinnor går nerför en gata.
En liten flicka som bär vit jacka sätter sig på trottoaren.
En tjurterrier terroriserar ett gammalt däck i sanden.
Ungefär 5 år gammal pojke, allt i svart, går på krusad strand.
En ung pojke lutar sig mot en stolpe med randig flagga.
En flicka cyklar i en korsning.
En svart hund jagar en boll i gräset.
Människor i rummet verkar arbeta på ett projekt men just nu äta och dricka.
Två unga män som arbetar i en trädgård.
En man i vit skjorta läser tidningen bredvid en man som bär mörka solglasögon.
Flera personer står runt i grupper bakom ett bord med bananer.
En ung pojke som hoppar på en studsmatta utanför ett hus.
En man som står på en bro under en kran.
En man i regnrock står i en torrdocka bredvid ett skepp.
En man med rött skägg kör en vagn längs en trottoar.
I ett gathörn står en man nära en hög med sopor sorterade för återvinning.
En kvinna som tittar på en mobiltelefon medan hon står på en trottoar.
En ung kvinna samtalar på sin mobiltelefon medan hon sitter på cementtrappor.
Två barn med björnseder sitter på trottoaren.
En kvinna som bär en lång svart läderrock och knäna höga svarta stövlar, med en stor blommig tryckblöja, köpa en tidning.
En blond kvinna bär en bricka med fyra små vita koppar.
Två damer med blont hår i jackor som går framför en stor byggnad.
Grupp av människor runt ett runda bord stapla spelkort.
En person i en stor svart hatt äter en skål nudlar med ätpinnar.
Tre personer står utanför ett varuhus.
En man som sitter på golvet bredvid en kvast en hink.
En svart man som bär en dunjacka med armarna utspridda och håller i en rosa kam.
Ett äldre par går nerför kvarteret under kvällstimmen.
Kvinnan i solbränd jacka står utanför och tittar upp.
En kvinna i turkos och brun rutig jacka som står på en gata.
En pojke i blå skjorta har ögonbindel och håller i en pinne.
En äldre djärv man med skägg i den ljusa skjortan sitter och röker på gatan.
En man som går genom en folkmassa på en stadsgata.
En man med solbränd jacka går in i Le Mignon på eftermiddagen.
En kvinna i svart går in i en tunnelbana under natten.
En man pekar på en projicerad bild av en Firefox-sida på en konferens.
Tre män målar en metallvägg vit.
Flera män sitter vid ett träbord på höger sida av gatan.
En flicka fixar sitt örhänge på sidan av en upptagen, bred trottoar.
En svart man sitter i sin stol och stirrar ut i fjärran.
En man i vit skjorta som sitter och övar ett musikinstrument.
En blond tjej som går och pratar på en mobiltelefon medan hon håller i en rosa plånbok.
En grupp människor samlas på gatan.
En konstnär i en grå t-shirt ristar på sin vita serpentinformade skulptur.
En kvinna i jeans går nerför gatan.
Fyra musiker spelar musik i en grupp på trottoaren.
En man i orange skjorta som går på en stig.
Människor som sitter vid bord med turkosa och vita paraplyer med utsikt över havet och stranden.
En man på en dammig båt som håller ett fiskespö.
Utomhus går tre kvinnor mot kameran när en av dem trycker på en barnvagn.
Turistfru upprörd med make som inte kan sminka sitt sinne.
En kvinna, som bär grå rock, lägger kläder i en tvättmaskin på en tvättomat.
Mannen ramlade precis av sin cykel
En asiatisk man som bär jeans och en blå knapp upp skjorta med en vit krage ligger på en parkbänk som håller en ljusfärgad jacka.
En tidig morgon rusningstid mitt i staden.
En gymnast ses trotsa gravitationen när hon utför ett imponerande drag flera meter ovanför de parallella barerna.
Ett litet barn bär en blå randig skjorta.
En manlig fotbollsspelare försöker leda bollen förbi målvakten för att göra mål.
En stor modern teater är upplyst på natten.
En ung dam som poserar med stolthet för en plats hon är stolt över.
Ett ungt barn som ler mot kameran medan hon står i trädgården.
En utsikt över byggnader och människor som går tvärs över gatorna i Times Square i New York.
Gamlingen gör något i sin verkstad.
Två äldre människor i bruna rockar står utanför och pratar med varandra.
Besättningen städade bort isen och snön från trappan.
Asiatiska turister stannar framför ett stort träd och beundrar dess rötter.
Tre äldre män är i en databutik.
En man klädd i blå och röd dräkt hoppar över en liten våg.
Gamlingen använder en improviserad trasig hjulpipa för att transportera sina verktyg till jobbet.
En kvinna som står framför en byggnad när andra gör sin dag.
En liten flicka njuter av en diet Coca Cola i en trädgård.
Shier i luften efter ett litet hopp i hans körning på sluttningen.
En man sitter bredvid en kvinna som står.
En hane som bär gula byxor fångar luft när han snowboardar nerför ett tomt berg.
En grupp människor går på trottoaren, medan en man letar efter något.
En tårta med fem vanliga ljus och ett högt, gnistrande ljus ligger på ett bord framför två män.
En skadad bil står parkerad mittemot folk i en grå bil.
En kvinna sitter på en berggrund medan man tar en bild och den tredje tittar ner.
En medelålders man som poserar med en krabba
En pojke använder ett baseballträ i plast för att öva på att slå en boll från ett slagte.
En man med metallföremål fastnade vid honom.
En besättning filmar en scen för en film eller TV-show på en gata.
En demonstranter som bär en USA-skjorta har en skylt under en protest.
Två män hukar sig ner på golvet och tittar på fyra hundar som leker i en bur.
En kvinna sitter och läser på en tvättomat.
En grupp barn färglägger lakan med kritor medan de sitter ett bord.
Ett band är i en inspelningsstudio och väntar på att börja spela.
En man klädd som en brandman sitter ner.
En kvinna som bär ett svart plagg håller i en penna.
Protester med politiska tecken samlas kring en musikalisk händelse.
En leende man har en skylt som föreställer en regnbågsfärgad elefant.
En man som poserar med en "november kan inte komma snart nog" affisch.
En djuraffärsanställd visar en skjortlös kund de olika typer av fisk som finns.
En kvinna går nerför en trottoar kantad av körsbärsträd i blom.
Två barn svingar medan de står.
En brun hund som hoppar i en stenig bäck.
En man sitter framför en butik i skuggan.
Många skjortlösa män, som bär svarta huvor över hela ansiktet, går barfota i en lång rad med en enda fil.
Ung barfota kvinna skrattar i hängmatta.
En man bugar sig i bön över en mycket utsmyckad kista i en katedral.
Folk gör sin dag i storstaden.
En man i svarta byxor och en grön polotröja plockar upp skräp runt sin mans sjö.
En kvinna i en stad tittar bakom henne.
En ung kvinna i jeans och en grå tröja går över en tom gata.
Unga flickor som uppträder någon form av dans.
En kvinna som bär förkläde står utanför en affär och pratar med en cyklist.
Barnen i blått sjunger för en grupp människor.
En munk i sin röda dräkt håller ett paraply utanför ett tempel.
En man i brunfärgad jacka pratar med en kvinna i svart kjol.
En ung man vit en vit, knapp-up skjorta, kör en blå cykel.
Vissa professionella baseballspelare värms upp.
En brunhårig kvinna som sover på en soffa med huvudet på en hög kuddar.
En kvinna går nerför en gata på natten.
En stor hund leker med en liten hund i smutsen.
Två barn håller upp fredstecken och ler.
En man i neongröna kläder knuffar en grön kärra nerför gatan.
En ung kvinna sitter på trottoaren och ritar en byggnad
En New York Mets spelare går på ett grönt fält.
En asiatisk kvinna står längs en väg där 2 bussar har passerat hålla sina väskor.
En flyktartist som bär Converse High tops kämpar på ena foten när en publik tittar på.
En kvinna som bar en stor väska på huvudet när hon gick nerför gatan.
En man som joggar på en fin park joggingstig, omgiven av vårens lövverk och träd.
Runner lämnar startblocken för ett lopp.
En man i brunt knuffar ner en container på en trottoar.
En kvinna stannar för att titta på några bröllopsklänningar.
Fyra personer hoppar på en sanddyne en solig dag.
En publik som går förbi med flera åskådare tittar på en gatuartist.
Människor går genom lobbyn med fläckar av dagsljus och skugga reflektioner.
Två kvinnor går nerför gatan och håller parasoller.
En staty och träd i en plaza framför en byggnad med människor som går förbi.
En man i stor skara samtalar med sina vänner.
En svartklädd man går över gatan.
En grupp människor väntar i en tunnelbana.
Två kvinnor, en i rött och den andra i vitt, är ute på joggingtur.
Kvinnor klädda i exotiska kläder, stående på gatan.
En kvinna med röda blommor står vid ingången till en byggnad.
Två par balettdansare uppträder utomhus.
En svart man pratar på sin mobil och håller i en vintagekamera.
Surfaren rider en våg tillbaka mot stranden.
En man som bär en säck längs en vattensamling.
En ung kille som hoppar ner i vattnet.
Två solbadare i skumma blå baddräkter ligger på den graffititäckta trottoaren.
Här är en ung man som skateboardar upp på sidan av en skate grop.
En man i en guldsmed sitter medan en annan man inspekterar sin sko.
Solen går ner när en man cyklar.
En kvinna klädd i vit skjorta, korta shorts och en fedora, går bort från kameran.
En man i gul skjorta skiner om ett tak.
En asiatisk man i traditionella kläder låter ett stort horn i ett behagligt bergslandskap.
En man i en baklänges hatt står i en Best Buy-butik.
En pojke njuter av att äta pizza i en tallrik.
Mannen går längs sidan av ett svart järnstängsel.
En medelålders vandrande man som bär glasögon och grå kostym täcker munnen med bilar som springer i bakgrunden.
En äldre man som tittar på en tidning när han korsar en gata.
Två män låter sina hundar leka tillsammans på gatan.
En man i röd skjorta och svarta byxor på stranden.
Två män som håller spadar står runt jord och träd.
En man spelar en xylofon.
Detta är en gatuscen med en hel del bilar och människor som går runt i olika riktningar.
Gymnast klädd i rött och svart poserar med åskådare i bakgrunden.
En kvinna som bär lila och bär en väska går ut genom en dörr.
Två kvinnor som pratar framför en gammal byggnad.
En cirkel av män i svart håller fjäderklädda hattar och står bakom ett rött tecken.
Väntar på tunnelbanan efter en lång arbetsdag.
En person sitter på en kulle med träd i förgrunden och målar en lugn bild av en sjö.
2 män som håller en skylt framför ett metallstängsel.
En cyklist verkar reparera en cykel som vänds upp och ner på trottoaren.
En film med två personer som sitter vid ett bord.
En vit man i svart kostym korsar en livlig gata.
En dam spelar gitarr och sjunger in i en mikrofon.
Två kvinnor i tajta jeans går nerför en gata, en med en shoppingväska.
Damen bär någon form av sko går.
Två japanska kvinnor i traditionell dräkt går genom ett trångt torg, en med väskor och en med käpp.
En bilist passerar förbi och en grupp människor sitter på en bänk.
Kvinnan i den gula jackan och bär en blå hatt verkar titta på något.
Tre vuxna och tre barn står eller hukar runt ett barns lila cykel.
En pojke i gul fotbollsuniform står på fotbollsplanen.
En pojke sitter vid vattnet och försöker mata en svan.
Människor klädda i traditionella japanska klädesplagg går i en procession genom en innergård belagd med marksten.
Två kvinnor i kimonos står tillsammans leende.
En kvinna med svart jacka och svart handväska som går nerför trottoaren medan hon tittar på sin mobiltelefon.
Orange och vit riskkottar vilar på gatuplattor.
En man i kostym blickar upp mot himlen medan han är runt hästar.
En kvinna som tvättar sin minibuss på en självservice biltvätt
En man som bär solglasögon, jeans och en svart skinnjacka hoppar i luften med armarna och benen isär.
Folk går upp och ner på den livliga stadsgatan.
En kvinna och hennes helgon bernard hund sitter på en bänk i parken en solig dag
En man i renässanskläder sitter på en tegelvägg.
En man i orange skjorta säljer bratwurst för en euro till en gammal man i blå skjorta.
Tjejen i en klarröd skjorta lyssnar på öronknoppar.
En man med en bollmössa pratar med en dam med händerna vikta över bröstet.
En man i isbjörnsdräkt står med ett tecken i protest.
Män och kvinnor hoppar och tar tag i varandra på offentlig plats.
Kvinnan i mörk skjorta står ensam framför en gul bil.
Kvinnan och flickan sitter i den bruna läderstolen.
Grupp av unga människor som spelar trummor medan en publik tittar.
En fluffig hund bär ett svart koppel i munnen.
En man som bär vita shorts rider en vattenskoterbil.
En man i svart jacka står mellan två träd och håller upp en skylt.
En ung man är i en affär som säljer korv och vin.
Fyra kvinnor med väskor på axlarna, som gick nerför gatan.
En man som sitter på avsatsen och läser tidningen.
En blond kvinna med kort hår som klipper en torsdagskväll.
En gråhårig kvinna som sitter på en röd bänk och håller en käpp.
En stor grupp äldre människor sitter runt olika utomhusbord.
Två äldre herrar i svarta shorts, som går på stranden.
Två asiatiska honor poserar för en bild medan en man verkar bära sina väskor.
Cheerleaders och idrottare poserar med maskot för ett foto.
Tre barn har vita och svarta ballerina dans i ett gym.
En brunett kvinna med en solbränd jacka som sträcker sig in i handväskan.
En ung dam som bär en vit klänning med en blomma i håret och ler mot kameran.
En kvinna och en man som sitter utanför.
En grupp människor som lyssnar på en man talar från en monter som heter "Teva Neuroscience".
Många människor samlas för att få gratis råd och information.
En tjej i röd skjorta och sönderrivna jeans springer fingrarna genom hennes blonda hår när hon ser framför sig.
En kvinna klädd i mörka färger som knuffar någon i rullstol.
En skara människor, några med skyltar, går längs en bred stig i en stads park.
En gammal man med en blå skjorta sitter i rullstol vid sin syretank.
En grupp människor i hopfällbara stolar och rullstolar sitter ute i solen.
Två kvinnor i Saris arbetar tillsammans i en by.
Selena Gomez bär en cream tank topp tittar på staden efter att hon klivit av planet.
En kvinna står framför en nöjespark.
En man i en krageskjorta som pratar med en annan man i solglasögon.
En man i vit skjorta sitter och lyssnar på musik.
En kvinna i röd skjorta och några jeans ser ut som hon grälar med en man i rött och en stor väska.
Två unga asiatiska kvinnor köper mat från ett japanskt livsmedelsföretag.
En kvinna i rosa skjorta tar ett foto av en fisk i ett stort akvarium.
En man med tröjan över huvudet står på en stolpe.
Kunden höll påsen medan undersöka apelsiner medan andra marknadsbesökare undersökte produkter vid andra tabeller.
Ett barn som öppnar ett födelsedagskort på en fest.
Tre unga kvinnor lutar sig mot ett räcke över en gångväg.
En man på en grönsaksmarknad pekar på något.
En man med långt rött hår, en brun skjorta och rutiga byxor säljer frukt på en marknad.
En man och en kvinna med cyklar i en park.
En man som bär randig svart och vit skjorta går tvärs över vägen, längs andra.
En man står med en grupp åsnor på en gård.
En svarthårig kvinna bakom ett podi håller tal för en stor publik.
En man som läser en meny på en restaurang.
Det finns människor som står på olika lägenhet balkonger interagerar med varandra och människor på gatan.
Två kvinnor äter ute på en restaurang
En grupp musiker uppträder framför en liten publik i en udda byggnad.
En sjukvårdare tittar på en brandbil.
Två män och en kvinna står framför en teater.
En kvinna som gör en smörgås i en affär.
En publik tittar upp på två personer som står på två balkonger i en byggnad.
En samling människor på gatan på natten.
En grupp människor samlades på natten utanför en tegelbyggnad.
Riotpolisen står framför en pöbelhop, inklusive en man i Batmandräkt.
Det står en man i dörren och framför ett träd.
En man som står ensam i en park.
En brandstege på sidan av en byggnad dominerar en urban scen i en gränd.
Två brandmän som skrattar.
Brandmän i full utrustning går upp för en stege.
En äldre kvinna talar på en mikrofon.
En man som bär en hatt med sitt ansikte upplyst står mitt i en cirkel av människor.
Två män spelar sina instrument medan en tredje sjunger.
En skäggig ung man i t-shirt och jeans läser en bok på ett utomhuscafé
Mannen i vitt pratar med kvinnorna vid bänken.
Fyra personers silhuett bär ett föremål uppför en kulle.
En man i skinnjacka och hatt som tittar ut i fjärran.
Det här är en vacker kväll med floden och solnedgången.
En kvinna står på ett gathörn.
En kvinna jobbar på en bar framför en neonskylt.
Tre yngre kvinnor sitter utanför och pratar.
En man som bär en blå skjorta driver en bankomat i ett rum med en bild av Fidel Castro hängande på väggen.
En ung kvinna, som bär en Carnegie Mellon-tröja, lyssnar på sina hörlurar.
En överviktig man i en blå och svart huva i tröja arbetar på en bärbar dator utomhus.
En man drar en tränare med två Geisha ombord.
Två män, en ung och en medelålders, arbetar på en liten dator med en skruvmejsel.
Ett poliskontor använder en cykel för att slutföra sina plikter.
Ett barn som sover med en nallebjörn och en filt.
En tjej som ligger ner i en bastu med bara en handduk på ser avslappnad ut.
Flera kvinnor i vit t-shirt bär varm rosa kort peruker står utanför i en stad.
En brud och en man i smoking på trappan.
Mannen i en långärmad svart skjorta, verkar vara engagerad i dans, framför en blå skylt som innebär information om specifika platser.
Tri-nivå byggnad med människor som står på varje nivå balkong som folk tittar på underifrån.
En man i en jacka lyfter armen omgiven av människor som är böjda eller huk.
En kvinna i lång klänning hänger kläder på en klädstreck.
Många möbler staplade ovanpå varandra.
En ensam vandrare som går på smuts med snöig fjällbakgrund.
En man med galna ögon i en fedora har sin gitarr tittat på.
En kille i svart läderjacka som riktar en ficklampa mot sig själv.
En man som interagerar med sin dotter på ett köpcentrum.
En gentleman i jeans och en svart tröja talar ivrigt på en mobiltelefon.
En tjej med en knapp ner skjorta med blont och rosa hår går.
En grupp människor som rider på en fullsatt buss.
En liten grupp människor står framför butiken och pratar om att hålla i en "Bönare Booth" lila skylt.
Människor i främst affärskläder skyndar sig längs en trottoar i staden.
Två män med målade ansikten ser ut som clowner en sjunger och den andra spelar en liten gitarr.
En liten flicka med ljusrosa byxor sticker lekfullt sitt ansikte i en tramption på en lekplats.
En ung flicka i rosa skjorta, blå jeans och sneakers som pratar in i ett objekt i en park.
En familj äter och tittar på TV.
Kvinnor klädda i en gul rock med en hane med ryggsäck på ryggen hugging mycket nära.
Studenter i en klass tar examen.
En kvinna i rosa och gul klänning går förbi en hög med däck och en gul grå randig byggnad.
Kvinna och man med käpp klättra trappor från tunnelbanestationen.
En man lutar sig mot en telefonautomat medan han läser en tidning.
En försäljare går nerför gatan och säljer sockervadd.
Det är tre killar som går längs trottoaren, den som är framför, jonglerar.
En man säljer dekaler på gatan.
En man och en kvinna på scen med en mimare.
En tjej i svart jacka som pratar på en mobiltelefon.
En liten pojke tar en bild med en digitalkamera.
En rad som väntar på att få komma in i en film
En man i svart bär shorts och solglasögon hoppar från en sten till en annan.
Snygg blond tjej som gör ett väldigt fult ansikte.
Två skyltdockor är i fönstret i en stängd butik.
Den här kvinnan och mannen har ett samtal.
En blond kvinna med blå skjorta går nerför gatan medan hon håller i sin mobil.
En man och en kvinna som står på ett berg har utsikt över det.
En man står vid två fordon med tre uppblåsbara amerikanska flagga designade fladdermöss lutade mot honom i en triangelform.
En man som säljer blommor, cigaretter och godis på gatan.
Två stövlar är på två skidor som rör sig väldigt snabbt.
En man som rider häst och leder andra hästar genom vacker natur.
En rad sadlade hästar går nerför gatan förbi en bil som har sin huva och stam öppen.
En röd spårvagn är på gatan.
Två personer promenerar framför en vietnamesisk restaurang som har graffiti målat på den.
En man och en kvinna som går hand i hand förbi en sportaffisch.
En ung man i en blå t-shirt går förbi en gränd medan han pratar på mobilen.
En man läser en tidning nära en gata full av fotgängare.
En man som bär på en väska håller handen mot huvudet och tittar uppåt.
Sex personer står vid räcket vid El Tambor.
En liten flicka i blå blomklänning och svarta stövlar som går på trottoaren.
Studenten tillbringar sina raster utomhus och njuter av varandras sällskap.
En kvinna och en flicka sitter under ett träd.
Två kvinnor i hatt går nerför gatan.
En man som sträcker på bålen i en motionsanläggning utomhus.
Man rider på en surfbräda på en våg.
Två skidåkare står på sidan av en snöig bergssluttning.
En gentleman med en grön jacka som tittar på en taggad vägg.
En ung man håller i en mikrofon med färgglatt ljus runt sig.
En man som fotograferar en stor betongvägg.
En grupp människor är på en nöjespark.
En man avfyrar ett spjut med en atyl-atyl.
En man i brun krage i skjorta stirrar ut i fjärran i en park.
En svart kvinna går till jobbet.
En ung pojke står på en gata med en påse runt halsen.
Män som för ett samtal nära en strand.
En man i blå jeans och en vit t-shirt som spelar saxofon
Arbetare under en motorväg som manipulerar ett metalltäcke på vägarbeten.
En kvinna som bär gult är ute under en hydda som ännu inte är helt byggd.
En pojke som tittar in i kameran och ett hus som byggs i bakgrunden.
En kvinna ler, håller en bok framför en folkmassa tittar på henne, i ett bibliotek
Minst tolv killar som bygger en byggnad, en del hjälper varandra.
En kvinna i jacka och pärlor på en boksignering.
En rad motorcyklar framför en affär.
En man som sitter bredvid en motorcykel på sidan av en gata.
En kvinna lutar sig mot en vägg med sin sko av.
En kvinna och två andra sitter i närheten en dekorativ vattenfontän.
En kvinna vid namn Victoria Leak sitter bakom sitt skrivbord på sitt kontor.
En kvinna klädd i vitt går förbi en byggnad som har en affisch på displayen.
Två vakter sitter nära en ingång.
Tre små blonda pojkar samlas vid basen av ett träd nära några gamla maskiner.
Folk hänger på räckena som gränsar till en gata.
Den asiatiske mannen får sin bild tagen med en motorcykel av en annan man.
En asiatisk man uppträder med ansiktsfärg på.
Två män är på väg att kliva av ett tåg.
En man med hatt är ute och annonserar en tatueringsaffär.
En skäggig man som bär målarmössa spelar xylofon på en livlig gångväg.
Ett skolband utspelat för andeveckan.
En ung dam som bär vinterjacka och gör sig redo att knäppa ett foto.
En livlig stadsgata på natten.
Flera människor sitter på en vägg täckt av graffiti.
En barfota man som sitter på en avsats vid en trottoar.
En person i röd hatt, slipsfärgad lila skjorta och svarta byxor står på en gångväg.
En man i grön tröja som springer.
Två smala svarta män sitter vid sidan av gångvägen, med varor att sälja.
En gammal dam och hennes barnbarn jobbar i en närbutik.
En asiatisk man i orange jacka bär en hög hög med lådor.
En man kör en kundvagn full av matvaror.
En man i solbränd jacka och blå jeans cyklar.
En uppsättning skådespelare och skådespelerskor utför en show.
En hona i en blå jacka som äter medan hon sitter på gräs.
Två kvinnor med paraplyer stående på en tågplattform.
En man och en kvinna äter lunch medan en kvinna i rött använder sin mobiltelefon.
Ett par som båda bär glasögon går och håller varandra i handen.
En kvinna med ett vitt huvudskydd rider en cykel på trottoaren i en stad.
Tjejen på en cykel går nerför en gata.
En kvinna med brun väska fäster en rosa och gul bukett på sin cykel.
Ett par bär påsar utanför.
En man håller upp ett tecken som lyder "Jobs with Justice".
En äldre kvinna tittar på en påse frukt medan andra tittar på.
En man och en kvinna som står mot en vit vägg och tar en bild med skuggor mot väggen.
En ung flicka läser en bok mitt i en stor röra av kläder.
En vit man och kvinna pratar, medan en svart man tittar på dem.
En liten flicka sveper utomhus.
Damen som håller en vit hatt går på trottoaren med sina två vänner.
Två barn, en av dem spelar trumpet för dricks
En äldre kvinna i en blå rock är på väg att prova ett prov av en röd vätska.
En clown gör publiken glad.
Ett par hemlösa människor rotar igenom en väska som innehåller saker som får dem att skratta.
Ett punkband spelar på scenen.
Människor i ett tält serverar och väljer mat och dryck.
Folk springer i ett lopp, två av dem bär färgglada indiska huvudbonader.
En kvinna som står på gräs, håller jackor och en klänning.
En man spelar trumpet inför en folkskara
En grupp barn samlas på stranden och pratar om vad de ser.
En elev observerar celler under mikroskop.
En man i gul rock, röd slips och clownnäsa pratar med en annan man på gatan.
Den unga flickan kom förberedd för regn.
En kvinna med lila paraply stirrar i fjärran.
Passerseglare som håller parasoller handlar grönsaker på en gatumarknad.
En man med dreadlocks och skägg pratar på sin mobil.
En kvinna och en man närmar sig.
Flera personer står på ett gathörn.
En utländsk marknad med en kvinna framför.
Det står kinesisk ung man och ung dam framför ett vitt bord med växter på sig.
Folk går på gatorna med paraplyer.
En man och hans hund går genom en fullsatt gata en regnig dag.
En man i en rutig kostym rock gester med sin hand.
Kvinnor i fina kläder har inget paraply.
En madrass lutar sig mot en telefonstolpe.
En man och en kvinna står mot varandra utanför framför en urna längre än dem.
Två kvinnor tittar från en bro på något.
Män arbetar på färgen på en sida av en gammal byggnad.
En ung flicka i rött är på en hopptur.
Två kvinnor kysser varandra på en cykel.
En liten lockig hårflicka som dricker ur en stor kopp.
Ett rött tält framför en tegelbyggnad betjänar förbipasserande på tegelvägen.
En stor skara av hundratals människor samlas på gatorna.
En man sparkas av en tjur när en rodeo clown springer upp.
Pappa och son bär matchande cowboykläder och tittar på rodeo.
En stor grupp människor samlas i en stor stad.
Det är folk som samlas utanför med flaggor.
Två personer i solglasögon pratar medan de sitter framför en stor gräsyta.
En man och en kvinna som sitter nära gatan.
Tre män har roligt när de använder den berömda vattencykeln.
Två personer klädda i gorilladräkter går längs en trottoar.
En stor grupp människor, några håller röda skyltar, nära ett gäng byggnader.
Folk som står vid startlinjen för ett lopp.
En man i svart skjorta går nerför gatan och erbjuder ett glas vin till en kvinna.
En kvinna med långt blont hår i en vit tank övredel håller upp armen.
En massa människor fyller gatan framför en McDonald's.
Tonårstjejen vill hjälpa till med smutsjobbet.
Folk går på gatan och konfetti faller på dem.
En grupp unga flickor som går nerför en gata.
En ung kvinna i jeans och en röd tanktopp sitter på en veranda med en ung man i halsband och shorts.
En kvinna i en röd topp som släpper Mardi Gras pärlor från sitt sovrumsfönster.
Två kvinnor i kavajer och jeans går genom en park och pratar tydligen.
Protesterande ungdomar koppla av i tunnelbaneparken, observerats av beväpnad polis.
Två honor, den ena i en rosa topp den andra i vitt, går nerför en gata
Brunett flicka ger förbryllad look samtidigt som bär en handväska.
En grupp trendiga ungdomar står utanför.
En kvinna med orange hår som sitter bakom ett bord med Tye-färgade t-shirts på sig.
En grupp kvinnor i stora hattar står vid ett bord.
En cyklist i blått parkerad inne i en träbyggnad.
En person i en folkmassa som tar en bild av människor på en scen.
En man som håller ett barn med ett barn på ryggen.
En man och en kvinna håller ihop, och en ung pojke och ett barn.
Två män som sitter bredvid varandra tittar åt olika håll.
Tre män sitter och en står och pratar med varandra.
En man i en bänk tittar på en annan man som sover.
En kvinna som bär glasögon håller en kamera i ansiktet.
En flicka i vita stövlar som håller i ett paraply.
En medelålders man i vit rock talar in i en mikrofon.
En kvinna i vit klänning går genom stranden en vacker dag.
En manlig ung man i svarta kläder bär en ryggsäck med en protestskylt i sig.
Man i jeans, knäpp upp skjortan, och bär glasögon läser en bok.
Ett barn med orange ryggsäck bär ett grönt fågelhus.
Mannen i den gula skjortan spelar musik på trottoaren.
Tre kvinnor med svarta kjolar möter en träddunge med lila blommor.
Ett par går förbi körsbärsblomträd.
En grupp människor står på stranden medan andra människor är i vattnet.
En man och kvinna boxas i en park.
En man och en kvinna står tillsammans när honan har en bit mediautrustning i handen.
Fyra unga flickor poserar för en bild.
En stor grupp människor samlas utanför en mycket upptagen gata.
Två kvinnor delar sockervadd på ett livligt stengator.
En man i blå skjorta följer en annan man som bär en blå och svart väska.
En tatuerad man får kroppsslag i en boxningsmatch.
En man har utsikt över en inredningsarkitekt på sitt hem.
En blond kvinna med en mörkblå tanktopp håller i en kamera.
En kvinna i solbränna lagar mat.
En mörkhårig man som röker en cigarett utanför.
En man i blå skjorta pratar med två män i orange och gul arbetsväst.
En kvinna som häller upp en kopp te.
En familj njuter av drinkar på däck med sin lilla pojke.
Två kvinnor handlar i en asiatisk närbutik.
En man sträcker ut armarna framför en stor klippformation.
En liten flicka rider på en brun ponny på gården.
Två små pojkar går mot en cykel framför en gul vägg.
En fotografering med en kvinna på gatan i röd och vit klänning och svarta stövlar.
Asiatisk man på en cykel som bär roller som matta och en annan kille.
En pojke tittar igenom några brädor på någon utanför.
En ung man och en ung dam som omfamnar under en täckt gångväg.
Två små hundar springer genom gräset.
Folk handlar på en utomhusmarknad för mat och kläder.
En person som håller en käpp sover på en bänk utanför.
En leende äldre man med vitt skägg och en äldre kvinna ser ut ett tvättbart fönster.
Sex kvinnor klädda i rött, stående på scenen.
En ballerina i en svart leotard hoppar genom luften.
En gatufruktförsäljare som väntar på kunder.
En ung man sveper trottoaren med en röd, hanterad kvast.
En tjej i randig baddräkt hoppar ner i havet.
Man i röd boll lock grillar fisk på grill.
En kvinna i gult går utanför en byggnad.
Uppifrån-och-ned-vyn av en man som sitter på en bänk inuti med en stående man vänd mot honom.
Fyra tjejer är på balett.
En man med solglasögon och en stor hatt med fjädrar poserar för en bild.
Två honor äter glasstrutar.
En man med svarta kläder sveper steg med en kvast.
En man står i en bäck omgiven av stenar.
En pojke och en flicka klappar en ko genom ett stängsel.
En man i vit jacka tar en bild.
Två män i blå skjortor står i tältområdet.
En man står vid en gatuförsäljares bänk i en stad.
Ett par äter utanför vid ett bord och han pekar på något.
Stor hund rullar på ryggen i grönt gräs.
En man i rosa knappskjorta höjer armarna framför folkmassan.
En svart och vit hund hoppar över ett hinder.
En disk i en restaurang med Marugas tomatpajer och baksidan av en Coca-Cola sodafontän.
Två killar i gatukläder som håller på med marshalkonst.
Två vänner håller i varandra och ler samtidigt som de njuter av en musikfestival.
En kvinna håller sitt barn under en fest.
En liten pojke sitter på sin fars axlar med ballonger i röd kostym.
Två svarta män tittar på en basketmatch på TV.
En kvinna i fuchsia shorts och en behå topp hoppar i luften.
En flintskallig man går på en stig skuggad av träd.
Två äldre män använder tång för att hämta mat från en frukostbuffé.
En grupp människor utför en fotografering.
Två asiatiska kvinnor bär sandaler, långa sidendräkter och håller parasoller.
En japansk man i blå hatt sitter med sin banjo.
En äldre kvinna som bär en blomskjorta väntar tålmodigt på att tåget skall stanna.
En man drar två kvinnor nerför en stadsgata i en rickshaw.
En gammal man som tvättar stadens fönster tänder böcker.
En man med solglasögon har grönt på armen.
Två kvinnor sitter vid ett bord i en cafeterian med blå, gröna och gula stolar.
På en stormarknad köper folk sina matvaror.
En äldre man i en rutig skjorta syr på en Singer symaskin.
En kvinna i en fin tröja hand gör något kreativt.
Ett par asiatiska människor står utanför nära en "rökområde" skylt.
En del japaner njuter av fyrverkerier från en lokal gata.
Två barn som sover i baksätet på en bil
En kille springer nerför fältet och håller i en fotboll medan hans lagkamrat, en motståndare, och domaren springer bakom honom.
En man i vita byxor och vit, strippad skjorta, och en kvinna med en kort svart och vit klänning dansar på ett kakel dansgolv.
En kvinna på ett blomsterfält blåser på dem.
En kvinna som sitter ute och väver en lång bit rött, vitt och blått tyg.
En ung flicka i alla rosa kläder som går.
En kvinna som går längs en betongväg ovanför havet.
En gammal man håller upp ett tecken.
En man som bär en röd jacka går på styltor framför en grupp människor.
En grupp blonda unga kvinnor sitter utanför en Star Bucks.
En flicka i grön skjorta tar en noggrann titt på ett objekt.
En kvinna står i dörren till en gammal byggnad.
Hunden bär en rosa boll i munnen.
En stor amishfamilj som ser längre än till en trevlig vårdag
En liten flicka i en ljus rosa hatt och rosa kläder håller en glass kon efter att ha gjort en röra av glass i ansiktet.
Tre gatuartister som visar upp sina extraordinära instrument.
Poliser tittar på som åskådare njuta av en parad.
En man går förbi en stor tegelbyggnad som är målad med graffiti.
Tre personer, alla med handskar, använder en skottkärra för att göra gårdsarbete en solig dag.
Cooks jobbar i ett kök.
Ett vuxet par i ett afrikanskt land poserar på ett rent smutsfält med en leksaksbil som håller en plastflaska.
En man i färggrann kostym med trumpet.
Två män går förbi en färgstark butik när man beundrar något under paraplyet.
En kvinna gnuggar papper på ett kakark i ett kök.
Ett foto på ett par som går nerför gatan med kinesiska tecken skrivna på skyltningen.
Ett ungt barn med blont hår försöker sätta en mobiltelefon i munnen.
En man och kvinna står framför en annons på en vägg medan hon tittar på den, han tittar bort.
Fem personer målar utomhus på trottoaren med sprayburkar.
En man med blå hatt och blå jacka stående på trottoaren.
En man i kostym går bredvid en vägg.
Dam med grått hår med mobiltelefon och bär en shoppingväska framför en butik.
En vacker kvinna som kollar sina mobilmeddelanden när hon går på en plaza.
En man med brun rock och blå huvudduk knäböjer och tutar en gitarr.
En blond kvinna med röd skjorta och fotbollshatt ler.
En mor och far tar sin på liknande sätt klädda familj för en promenad i det offentliga området.
Mannen i jeansjackan tittar tvärs över gatan.
En man i jeans med röda skor cyklar nerför en gata förbi en tegelbyggnad.
Damen är grön håller i ett bindemedel.
En man i rutig skjorta röker en cigarett på en gata.
Två män och en kvinna utanför ett bostadsområde.
En brunett kvinna med en lei på huvudet som sticker ut tungan.
En kvinna ligger ner i gräset i en park.
En man i rosa skjorta syns dricka en öl.
Folk tittar på en tävling på stadens gator.
En man i färgglada kläder och hatt står i en folkmassa.
En gymnast med hjälp av en uppsättning parallella barer.
En man fäster färgade svampar på skjortan och jeansen.
En man böjer sig över med ett uppstoppat djur mellan benen.
Två unga damer i en bandgrupp med trumpinnar.
En kvinna med en trumma leende
Mannen med rakat huvud hänger upp tvätten på linjen.
En gammal man som tittar över en skulptur.
En kvinna i lila skjorta och rosa hade gått i en skara människor.
En man är klädd i lila och orange kläder för en händelse.
En kvinna klädd i en gyllene dräkt ser ut att vara på avstånd.
Man i puffig gul jacka på skidor på ett berg.
En grupp människor tävlar med en man klädd i drakdräkt.
En kvinna tar sitt barn på cykel.
En kvinna som går och bär en ljus rosa rock och kort, tight svart klänning.
En hund går utmed en röd tegelgata.
En svartklädd man sitter vid en lyktstolpe och röker en cigarett.
En kvinna som viftar med den mexikanska flaggan.
En kvinna ler mot ett barn i en barnvagn på en äng.
En skara människor som viftar med sina armar.
Folk ställer upp sig och gör sig redo för Flag Day i Frankrike.
En man i en grön hatt dozes när du rider på tåget.
Flera personer inklusive ett barn och en clown går mot en snöig trottoar
En grupp äldre kvinnor som sitter på en bänk med samma hattar.
En man i svart skjorta står upp och gör bubblor.
Tre personer sitter på sina bärbara datorer i ett kafé.
Två män klättrar upp för en stor sten.
En man som går på en grusväg.
En grupp på sju kvinnor står i en vattenförekomst.
En ung asiatisk man sitter bakom ett schackbräde och väntar på att den andra spelaren ska komma.
Barn tävlar i en potatissäckstävling vid en utomhusfest.
Tre personer gör armhävningar.
Män spelar olika musikinstrument i en park.
En man och en kvinna dansar.
Barn tittar upp på en bronsstaty av en häst och en soldat.
Grupp av människor, mogna och unga sitter bredvid grusvägen tittar över vägen.
En man i 30-årsåldern sitter på en trottoarkant, klädd i en pälsig grön kostym.
En flicka i rosa spelar trummor.
Två kvinnor står i snön och tittar mot ett torn med orange konformat ljus.
Någon med en cykel köper produkter.
En äldre man och kvinnor använder datorer i ett slags förråd.
En gymnast balanserar på en balansstråle.
En kvinnlig gymnast i en röd och blå leotard gör en backflip på balansbalken.
En kvinna håller handen mot ljuset när en man tittar på.
En man sätter upp eller tänder lampor.
Fotografer tar bilder på ett bröllop.
En man som tar en bild av flera personer, inklusive en man i en limegrön kostym.
En man spelar akustisk gitarr, medan en annan följer med honom på dragspelet.
En grupp turister som går runt på den vaticanska gården.
En gammal man spelar dragspel på trottoaren.
En blond kvinna håller sitt glas uppe i en bar.
En man som sitter vid sidan av havet och håller i en pipa.
En vuxen man kastar ett barn i luften på en strand medan ett annat barn tittar.
En blond kille i orange skjorta som leker med leksaker.
Två mopedentusiaster, varav en bär handväska, har ett samtal på trottoarkanten.
Folk går nerför en trottoar kantad av pastellfärgade byggnader.
En kvinna i en rutig skjorta nära en gata med tummen uppåt.
Tre barn tittar på männen som jobbar utanför fönstret.
En idrottsman som har glasögon som faller av sitt ansikte ligger i en sandlåda.
Någon sparkar en boll som är mångfärgad.
En gammal man med en påse chips sitter med en yngre man som håller i en drink.
En pojke med ett stort leende på gömt ansikte, på ett blomsterfält.
Två män går längs en väg i ett tropiskt område med en tämjd elefant.
En frisör i en salong tittar ut genom salongen.
En äldre man som sitter vid ett bord i en tom restaurang.
En man kastar pilen.
En vuxen man och två barn av asiatisk härkomst hoppar i vägen.
En man i röd skjorta som kastar en pil.
En svart hund är i gräset med en kvinna i jeans.
Två unga flickor med solglasögon sitter utanför.
En ung afrikansk kvinna stirrar på en kamera framför ett gäng lerkrukor.
En kvinna sitter på en parkbänk och äter glass.
En kvinna i gult, och en kvinna i orange, båda med handväskor, titta på vattnet i bakgrunden.
En blondhårig kvinna som kisar och bär en klargul skjorta.
Två unga kvinnor går, en lång, blond, modell-liknande är i en zebra stripe outfit, den andra kortare asiatiska i en vit chemise.
Två kvinnor i tank toppar och solglasögon går tillsammans.
En flintskallig man som står vid sidan av en t-shirt-display.
En liten pojke som jagar en svart kråka.
En ensam kvinna i röd skjorta stirrar uppåt med en man i glasögon som tittar mot henne, på avstånd.
En kvinna i solglasögon håller i ett paraply.
En kvinna leker dragkamp med sin svarta hund i ett brunt landskap omgivet av träd.
Två kvinnor går nerför gatan i staden och länkar samman vapen.
En kvinna i en blå rutig skjorta och solglasögon kliar sig i ansiktet när hon går nerför gatan.
Kvinna i hatt karusell på gatan med shopping väska i bärgning.
Tre personer spelar fotboll, en bär orange, två bär blått, varav en är mitt uppe i luften.
Två kvinnor går tillsammans.
En man i en svart grafisk t-shirt klädd i en vit handduk över den nedre delen av ansiktet.
En kvinna med kamera går längs en mans sida.
En arbetare är på en körsbärsplockare i en palm.
En skjortlös man hoppar med skateboard.
En flicka i solglasögon går förbi en röd bil.
Han äter maträtt och njuter av den.
En flicka går på en trottoar med hörlurar i öronen.
En man i gul och blå rock som ber en kvinna om hjälp.
En mycket rynkig kvinna som håller sina glasögon och går nerför en gata.
En uppsatt polis passerar en mc-förare.
Unga i blå jeans väntar på sin blinddejt i parken.
En kvinna på sin mobil går i en park.
En grupp människor sover på en buss medan en pojke skickar ett sms.
Ett nyhetsankare filmas i en butik.
En kvinna som står framför en stor tank på ett akvarium vänder sig om för att titta på fotografen.
En kvinna som står utanför en affär försöker stänga sitt paraply.
En kvinna och två män går på en uppsättning utomhustrappor bredvid en annons.
En kvinna i kostym med kondomer i håret.
Två personer bär blomkostymer och går nerför en gata.
En pojke tittar på en båt fylld med sand.
Två tonåringar, en man och en kvinna, bär sportuniformer som springer efter en boll.
Mannen i grå jacka sitter på bänken och läser en bok
Flera män bär röda mössor, en står skilt från de andra och tittar mot kameran.
Många människor går längs en trottoar.
En kvinna i röd rock korsar gatan med en flicka i röda byxor och en barnvagn.
En asiatisk man tillagar mat på en disk bredvid en katt.
En grupp äldre damer som står på ett gathörn i en urban miljö.
Folk som bär väskor går på en gata med en parkerad motorcykel.
Två skjortlösa män på en byggnad balkong pekar mot himlen och observerar något intressant.
En kvinna dansar bredvid en scen under en musikfestival.
En ung asiatisk flicka klappar ett djur av något slag och djuret lägger sig ner och njuter av det.
En hund hoppar i luften och fångar en frisbee i munnen.
En man sitter bredvid en staty av en annan man sittande, ser mycket lik varandra
En kvinna i solbränna som knuffar en barnvagn.
En gatumusiker sitter på en gata bredvid en didgeridoo och håller ett blått ägg-formade objekt.
Vänner och familj samlades utanför Papa Johns.
En kvinna stannar vid en korsning och väntar på signalen att börja gå.
En grupp medelålders människor rider en häst dragen vagn medan de är klädda i historiska dräkter.
En grupp coeds spelar fotboll medan de dricker.
Två män med ryggsäckar väntar.
En kvinna som hoppar som en man tittar på henne i luften.
Två unga kvinnor sitter i ett träd.
En arbetare med en vit hårdhatt är på botten av en yttre brandstege och kämpar för att arbeta med kanten av en stor gul skylt.
En man i kostym har precis gått över gatan.
En kvinna som står i en mörk dörröppning och väntar på att släppas in i byggnaden.
En hund följer en annan hund runt hörnet men ser tillbaka.
En ung flicka som flyger blå tights i flottan deltar i ett långt hopp, medan folk tittar på henne.
Tre personer samlas runt ett bord för drycker.
En individ skickar ut sin cykel i luften.
En pojke cyklar i en skatepark.
En pojke cyklar nerför gatan med en stor gul citronformad skylt medan en mängd människor väntar i kö på trottoaren.
En kvinna i en blå skjorta som griper en annan kvinnas rumpa.
En kvinna som sitter på trappan med mörkt hår och lägger handen på ansiktet.
Ett par står på en brygga vid vattnet och kramar.
En brud en brudgum får sin bild tagen på en swing uppsättning medan en ung man dricker en läsk och en pojke i en grön skjorta med en cykel tittar.
En ung flicka bär rosa rengöring stenar i vatten med en tandborste.
En kvinna som håller i en korg och bär en silverfärgad peruk med nya glasögon.
En kvinna och en flicka undersöker en målning.
En man i blå skjorta hjälper en man i röd skjorta fixa en trail bike
En dam som spelar musik på sin harpa.
En kvinna är uppklädd och försöker sälja sina varor som en ung kvinna ser på.
Två hinderare hoppar ett hinder på en bana.
Två barn som bär hatt hänger fast vid bambuträd.
Två män pratar medan en håller i en kyckling.
En äldre kvinna står på gatan och poserar i rök.
En asiatisk kvinna som bär jacka och håller i ett papper.
En man i en tröja håller i en lampa.
En man håller upp armen mot ljuset.
En dam står upp och hullar en lampa som är tänd.
Män förbereder en kanon framför ett slott.
En ung man spelar foosball med ett par andra människor.
En grupp på fyra personer samlas på en trottoar.
En man som bär en töljacka och håller i ett rosa paraply och går bredvid en kvinna i svart rock och går en hund.
En tonårsflicka som bär flanell hoppar på ett gräsfält nära en fotbollsplan.
En målning av en livlig gata vid Oxford Circus Station.
En arbetare med en hård hatt som arbetar på en rigg högt från marken.
Två barn kliver över toppen av stenar som skär en stig över den grunda floden.
En man och ett barn går över vatten med hjälp av stenar.
Flera ungdomar går över vattnet på en rad språngstenar.
Barn leker tillsammans i en översvämning nyligen.
En kvinna klädd som en magdansös går bakom tre personer som sitter på trappan.
Kvinnan sitter i skuggan med en tygfläkt.
Folk står utanför ingången till Fulton St Stations tunnelbana.
En man i mörka kläder som går på en transitstation.
Två stadsarbetare klädda är orange städar upp en brinnande röra på en stad gata och trottoarkanten.
De två mormor pratar med varandra.
Två äldre damer delar lunch på en bänk.
Två personer sitter nära ett träd och slappnar av.
Tre personer går över en stenbro på en sjö medan en hund simmar.
Två barn använder betongblock för att gå över vattnet.
Tre personer klädda i randig, rosa och grön skjorta ser på och samtalar med andra
En väntande lounge med passagerare som väntar runt på blå sittplatser.
Asiatisk brud och brudgum lämnar en kyrka med folkmassor som kastar konfetti på dem.
Två små flickor bär rosa klänningar och sandaler
En gata i en stad med bilar och byggnader.
En kvinna i rosa skjorta gör apelsinjuice på en restaurang.
En söt lockig flicka som sitter på en mans axlar.
Fyra tjejer spelar hopprep i orangea jackor.
Två barn bär orange väst och blå byxor, medan en tar en bild med en röd kamera.
En kvinna och två små flickor som leker med hulahoops.
En man sitter i en trehjuling med en skylt i ryggen som lyder "Din annons här!"
En man i en bandanna möter tjejer i blå skjortor.
Två unga kvinnor med brunt hår sitter på en trottoarkant.
En stor grupp individer samlas runt ett starkt ljus på natten.
En levande teatershow med fem skådespelare på scen som gör en koreograferad rutin.
Ballerina uppträder som en tjejråtta i en öppen park.
En man med en machete som hugger stora isblock.
Två flickor läste ur en bok tillsammans.
Tre män och en kvinna har bärbara datorer och står framför en projektionsskärm som verkar konversera.
En polis vakar medan många människor deltar i ett maraton.
En ung kvinna i en mörk tank topp och orange solglasögon spelar trummor.
Två gitarrister samtalar på scenen.
En man spelar gitarr framför ett stort tecken, med en annan man som spelar trummor bakom sig.
Ett band som spelar utomhus för en fördel i New York.
En kvinna med en blå rutig skjorta och en bandanna gör bröd.
En man stöter bort en klippa över vatten.
En man i rostfärgad hatt och brun skjorta som pratar in i en mikrofon.
Kvinnan i grön och vit randig mössa står nära graffiti.
En grupp kvinnor står på en marknad medan en del av dem bär korgar med grönsaker.
Två gamla kvinnor sitter på trottoarkanten bredvid blommor
Polisen fyller en gata fodrad med åskådare i röda kläder.
Ett band som uppträder på en utomhusscen.
Tre män spelar trummor och gitarr på scenen.
En staty av en kvinna med långt hår
Ett afroamerikanskt band spelar utomhus på en scen omgiven av träd.
En svart man i brun skjorta och hatt talar in i en mikrofon.
En man med lila bandanna är klädd i polisupploppsutrustning, inklusive en hjälm och en väst märkt "Polisen".
Många människor tittar på produkter till salu.
En pojke i gul skjorta springer i ett lopp
Tre personer går förbi en vägg med en tavla av en läkare som kollar ett hjärta på en "I heart NY"-affisch.
Asiatisk flicka spelar Jenga fruktar att bitarna kommer att falla över.
En fattig svart man har ett religiöst tecken medan han står utanför ett matstånd.
En man i röd skjorta och en man i blå jacka diskuterar och pekar på en plats på ett litet krukträd.
En liten flicka hänger på baksidan av en basketkorg.
En man som bär en grön skjorta och bruna byxor, verkar vara mycket spännande, hoppa i luften med händerna upphöjda.
Två asiska män använder sina färdigheter i träbearbetning.
Tre personer, två kvinnor och en man, samlas runt en grill utanför.
Två män rakar huvudet skalligt.
En man hukar sig över sina växter med olika växter och smuts i bakgrunden.
En flicka som bär cykelhjälm och glasögon tar en bild av några växter.
Kvinnan som bär scarfen väntar tyst på tåget.
En sångare i svart skjorta spelar i ett band.
En liten flicka i rosa kjol bredvid en pojke.
Två små flickor som leker tillsammans i sanden.
En man i bast och läderjacka som skriver i en liten anteckningsbok.
En långhårig kvinna sjunger in i en mikrofon.
En grupp äldre människor som spelar schack i ett mycket fattigt område.
Två äldre herrar spelar schack.
En man sitter mellan en orange käpp och en orange blomkruka med huvudet böjt.
En kvinna, som bär en rosa väska och ett vitt paraply, går nerför en tunnelbana.
En kvinna i en grön tröja som stirrar ner i vattnet från en bro.
En tjej i svart skjorta med blå jeans har ett silverhalsband.
En ung kvinna i svarta byxor står bredvid sin cykel och tar ett fotografi.
En asiatisk kvinna som går längs en upplyst stadsgata på natten medan hon pratar på sin mobiltelefon.
En kvinna i en hög bergskedja häller upp dryck från en kopp till en annan.
Mamma åker genom parken med grabben i bärgning.
Män som sitter på sidan av en tegelväg.
En smutsig man tar en tupplur på en offentlig bänk.
En person med blå hatt och byxor ligger ner med huvudet på en bit bagage.
En man lägger undan disken.
Två män som bär ryggsäckar går på motsatta sidor av gatan.
En kvinna väger något medan en man sitter ner.
En man tittar ut genom ett byggnadsfönster medan han står under en puertoricansk flagga.
En gatuförsäljare som sitter på en trottoar med ägg och levande kycklingar.
En grupp hundar fastbundna vid en stolpe en varm sommardag.
En man sjunger och spelar gitarr på scenen.
En musiker i en färgstark skjorta verkar utföra ett solo på en rutschkana gitarr vid en fullsatt utomhusmusikal händelse.
En mexikansk man rider på en kärra dragen av en åsna.
En pojke och ett barn som sover på gräset i solen.
Tre män äter lunch på en parkbänk.
En man i svart kostym spelar en brun gitarr.
En hund går nära en vattenförekomst.
Ett litet barn i gul jacka, rosa stövlar och en scarf går iväg genom en isig vinterpöl tillsammans med sin hund.
En grupp på fyra personer på tre skotrar stannade.
En person i röd kostym kör motorcykel.
En man är klädd i turban och en blå och brun morgonrock.
En kvinna med vit skjorta och jeans rider en motoriserad skoter.
En man sträcker sig samtidigt som han håller fast vid ett metallstängsel.
En man som har lite kul i Harlem under en av Halloweens högtider.
En skolvakt för att hjälpa barnen.
En gammal man som sitter på en buss och håller i en portfölj.
En blond kvinna i brun säljer räkor.
En gatuförsäljare lagar mat under en enda glödlampa på natten.
Kvinnan i hijab kör en scooter.
En tagghund biter en annan brun hund medan han ligger på en säng.
En kvinna som knuffar en barnvagn promenerar förbi en stor annons.
Två attraktiva kvinnor promenerar nerför en fullsatt tegelgata på natten.
En taxi med många människor runt gatan.
En ung asiatisk kvinna går förbi en blå vägg som säger "Post No Bills".
Flera människor korsar gatan vid en korsning.
En grupp ungdomar passerar några fordon och en graffiti utsmyckad vägg när de tar sig genom staden.
En kvinna i skuggorna med en rödhårig trasa runt halsen.
En kvinna som bär ett hjärtformat halsband och en blå skjorta är bredvid ett staket.
En grupp damer som ler för en bild.
En man med en cigarett lyssnar på en annan man i klädesplagg som håller en burk.
En attraktiv kvinna som går på en gata i en gul skjorta.
En fotograf i blå skjorta som röker mitt på gatan.
Sju tonåringar går genom en betesmark.
En man och en kvinna som står nära ett skrivbord medan en annan kvinna sitter vid skrivbordet och tittar genom ett mikroskop.
En grupp människor som står utanför en byggnad.
En man med blå jacka och glasögon sitter på en pall.
En man och en kvinna som har ett samtal och båda bär hattar.
En tatuerad kvinna med en grön klänning och gul ryggsäck som håller en vattenflaska går tvärs över gatan.
En ung man tittar och tänker samtidigt.
En man med långt svart hår som går nerför en gata i en asiatisk stad.
En person i en grön skjorta med ett färgglatt paraply.
En man som roar en kvinna och flicka på benförlängningar med en topphatt.
En man låser upp en blå garagedörr.
En person sitter på en avsats vid en flod i en stad.
Två män arbetar med en stege i Amsterdam.
En man med grå jacka och grått hår tittar på någons sko.
Precision är nyckeln när vakten kastar sin pistol i luften redo att fånga den.
En australiensisk fårhund sitter på en träbrygga, bunden till en vit segelbåt.
Två ballerinadansare uppträder på en scen.
En kvinna i en blå tröja, som håller i en kamera, hoppar i en park.
Två brunetthonor som bär solglasögon utomhus.
En man och två barn, ett barn sitter på en kudde, stirrar ut på ett akvarium fullt av tropiska fiskar.
En man i blå shorts boxas en annan man i svarta shorts.
Folk står i kö framför en butik och annonserar öl, is, vin och tobak.
En man med skägg pratar på mobilen och står bredvid någon som ligger på gatan.
Tre uniformerade arbetare städar utomhusfönstren på en restaurang.
En man i svart skjorta är på en skateboardpark som håller sin skateboard.
Två män spelar catch med en fotboll i en gräsbevuxen fält på en solig dag.
Olika människor korsar gatan av en spritbutik och Thai House.
Två män med gula västar hänger med slutna ögon i två cykelrickshaws.
En kvinna som visar en ung dam saker.
En man och en ung pojke som bär randiga skjortor går på en grusväg längs vattnet.
Två poliser går nerför stranden.
En dam går över en väg med ett paraply för att skugga henne från solen.
En man lutar sig mot en vägg med skorna av.
Man med skålklippt och grå skjorta fotograferad bakifrån på en tunnelbana.
En serviceman som bär en hård hatt sänks under en trottoar.
En kvinna i en vit tank topp sitter nät till vatten med en duk i knät.
En grupp byggnadsarbetare kikar ut i staden.
Ett par står utanför en tysk restaurang och undersöker menyn.
En grupp människor njuter av ett enat kall.
En man är klädd i poliskläder med hjälm och sköld.
Familjemedlemmar njuter av en vacker solig dag i parken.
En kvinna med blont hår, bär blå jeans, går förbi en musikbutik och lång, beige byggnad som har höga glasdörrar.
En ung pojke i röd skjorta står på en pall i ett badkar.
En man böjs över av en gammal stenmur, tittar in i sin ryggsäck.
Fyra kvinnor poserar för en bild.
En kvinna med brunt lockigt hår, med solglasögon, stående i en publik.
En kvinna som ligger på asfalt mitt i en livlig park.
Pojke med vitt pulver och blå skrift i ansiktet
En kvinna med röd rock med svart huvudduk står mot en vägg.
En äldre afrikanamerikansk man griper tag i något som går längs gatan.
En grupp flickor i svarta och vita fläckiga kjolar korsar en gata.
En man håller två flippers medan han står framför en båt.
En hemlös medelålders man som håller en läskkopp tittar på två personer som gått förbi.
Sidewalk konstnär koppla av på stoop efter en hård dag på kontoret.
En grupp människor stirrar uppåt, en del verkar vara i chock.
En person i vit skjorta som står framför en byggnad med mycket glas.
En mor och dotter som går på en gata.
En man i björndräkt, som håller kostymens huvud i handen, står bakom en folkmassa.
En dansande poledans mitt på gatan utanför BUA.
En person som sitter i en båge fäst vid en stolpe på natten.
Många människor samlades i en park.
En hona akrobat är suspenderad i luften medan du gör en slående pose
Den unga damen dekorerar sig själv för Halloween.
Patroner väntar vid och i närheten en korsning i ett främmande land.
En skäggig man använder verktyg för att rista ett träföremål.
En del män och en del kvinnor står utanför medan de bär färggranna kläder.
En man som sitter i en stol framför en vägg av bilder.
En skäggig man, som använder en trästolpe, rör skålliknande föremål runt i en stor metalllåda fylld med vatten.
Två män klättrar.
En kvinna skakar hand med en annan kvinna, medan de står under ett tecken för en protest de för.
Två japanska kvinnor håller kvastar och går på en trottoar.
En man med orange skjorta serverar snökoner från en glassvagn.
Flickor förbereder mat att äta.
En man bredvid en cykel med en flagga fäst för att få uppmärksamhet av andra runt honom.
En flicka firar sin examen utanför.
En man i grå skjorta går bredvid en betongvägg.
En man som väntar på bussen.
Tre barn är i stora uppblåsbara bubblor som flyter ovanpå en pool.
En liten flicka i blommig rosa kläder gråter.
Polisen i upploppsdräkt går nerför en gata.
En manlig löpare tittar på en annan när de tävlar.
En kvinna sitter på några steg och slappnar av med slutna ögon.
En man på en cykel hoppar från en ramp.
En BMX-cykelcykel i luften, efter ett hopp från en byggd gruskulle i en skogsmiljö.
En kvinna och en man dansar på gräs.
En man i en hatt stirrar framåt med folk bakom sig och bredvid honom gör samma sak.
Två kvinnor paddlar kajak på en stor flod.
En boxare i vita shorts får ett slag i ansiktet på boxaren i de blå shortsen.
En tjej som är inblandad i en omgång "Människo Bowling".
En man i svart jacka går sin lilla hund i ett pittoreskt område.
Arbetare i ett företag skär plast för en väntande kund.
En pojke står i gräset och viftar med sin nations flagga.
Flickor dansar bakom en man i vit morgonrock och turban.
En man framför en sjö som städar fisk i randig skjorta.
En kvinna som håller i en bricka med spritshots.
En ung gentleman med brunt hår, med solglasögon ovanpå huvudet, njuter av en uppfriskande drink när han går igenom en meny.
Pojke som kikar i en tjejs kläder på sin tatuering.
Många människor väntar i långa köer för att få köpa biljetter.
Taxibilarna kör nerför ravinen i regnet.
En fullsatt trottoar med människor på den skild från gatan av metallbarriärer.
En man lutar sig mot trädet och spelar klarinett medan han spelar in sig själv med en videokamera.
En gatuförsäljare med vita byxor och svart t-shirt står nära sin vagn med kalla drycker.
En man i röd skjorta gör något med ett cykeldäck.
En man i röd skjorta tittar på några saker på marken.
En ung man som lutar sig mot ett gatuljus som en buss med en staty av Liberty skylt kör förbi.
Två män ser tankfullt ut från sidan av en bro.
En kvinna som bär en tanktopp håller i ett blått paraply och knäböjer bredvid bagaget.
En grupp människor i ett främmande land några bär paket, komma promenader, några stående.
En fullsatt gata full av asiatiska människor.
Ett litet barn sitter utomhus på en grön och vit handduk och barnet ler mot någon till höger.
Grupp av människor på ett torg på solig dag
Två äldre människor, en man och en kvinna, sitter på en bänk med en stadsbild i bakgrunden.
Det här är bilden av en kvinna i en blommig klänning, som tonar något i en hink.
Två unga flickor är placerade bakom ett bord täckt av olika leksaker och miniatyrer.
En gammal man grillar mat på en bakgård.
En kvinna med rött hår står bakom ett staket med sin kamera, längs sidan andra människor.
En manlig artist handlar en historia för små barn
En kvinna i en orange halsduk har en vit mobiltelefon.
En person reparerar en cykel medan fyra personer tittar i en urban miljö.
En asiatisk kvinna bär en svart examen keps och klänning leende på en gräsmatta.
Två män spelar schack på en grön låda bord.
En pojke sitter på en röd stol och tittar igenom en bok med gitarr och förstärkare bredvid sig.
Två kvinnor går genom en urban miljö med campingutrustning.
En man med grå hatt spelar fiol.
En ung kvinna i ceremoniella kläder som går med parasoll.
En ung man häller te från en vattenkokare i ett glas.
Mannen i röd jacka är ointresserad av parad.
En ung man sitter på gräset och lagar något slags sportnät.
Många små segelbåtar sitter vid en brygga.
Make och hustru på väg uppför kullen för att gå till badhålet.
En man i en fez håller ut en kopp på en torgplats.
En afroamerikansk man står på gatan med en skål bananer på huvudet.
Två män spelar fotboll på vad som ser ut som en dyster dag.
Ett bi ovanpå en blomma
Vissa människor går och andra sitter vid ett gathörn.
En ung far i orange byggnadsväst har en ung son på axlarna som bär en matchande väst.
En kvinna och barn som svänger på en däckssväng.
En vacker dag för cyklar och motorcyklar, och att ha en bar-b-q med familj och vänner.
En man som sitter vid ett bord och röker.
En man och en kvinna jobbar hårt för att städa upp efter en lång dag.
En man skrotar färg från ett fönster.
En skrattande kvinna håller en rosa stjärnformad lampa mot huvudet på en skuggad person i förgrunden.
Två barn med rakade huvuden, ett med en käpp, stående på gatan.
En kvinna i Vegas ser ut som en showbruddräkt i en blå och vit befjädrad huvudbonad rör sig framför en skara blåskjorta individer.
En man äter på gatan när han går.
En liten flicka svänger högt ovanför ett trästängsel på gungan.
Bald man i kockens tunika greppa tidningen med övertygelse.
Den vackra damen häller något i den andra behållaren.
Två personer kramas bredvid en grupp tonåringar.
En man i en blå jacka som sitter vid bordet och läser framför en restaurang.
Två barn sitter ner omgivna av olika typer av mat.
En ensam bicyklist rider förbi en utsmyckat dekorerad tvåvåningsbyggnad med många fönster.
En motorcykelförare hoppar i luften medan någon i bakgrunden tittar.
Mycket mörkhyad man ser tillbaka på kameran bakifrån buffé.
En man som gick förbi en sittande man på gatan.
En gammal man som bär bandanna och ett denimförkläde tittar på ett skåp i en verkstad.
Denna smuts cyklist njuter av loppet på racerbanan i Atlanta.
En kvinna som stirrar på kameran bakom solglasögon, håller i en väska och kaffekopp.
En flicka skateboard i röda skor på trottoaren
En skjortlös man med en blå skateboard utför ett trick.
En kvinna går förbi en byggnad märkt Fisher's Popcorn.
En ung man står nära sin cykel utanför en butik som heter, "Saras Old Fashioned Ice Cream."
En kvinna i svart tank topp och nyanser med en tatuering på armen.
En man i vit skjorta fixar däcket på en crimsoncykel.
En hund hoppar över en hög med stockar.
En kvinna i svart skjorta och vita skor som pratar i telefon.
En skjortlös man i en vit stol ser ut.
Folk går längs en gata under en stor skylt.
Den här pojken går nära en gata.
En ung flicka som spelar krocket och ler eftersom hon mår bra i sitt spel.
Folk äter vid borden framför en konstdeco-vägg.
En dam går ut ur en kort tunnel när en man förbereder sig för att gå in i den från motsatt sida.
Gamla människor som står i en cirkel på en fest
En man med en mörk jacka, skjorta och byxor, stående nära en grill med en hand som håller i handtaget på grillens lock.
Barn gör olika saker i bilden, äter och poserar.
Fyra kvinnor ror sig nerför bäcken i kanoter med bambustjälkar och halmtak på sidolinjen
En flickas hår flyter bakom henne när hon svänger
En kvinna i svarta jeans och en bikini kastar handen i luften medan hon är på stranden.
En man njuter av solen i en park.
En grupp trogna shoppare bär kylan medan man pekar på hans favoritaffär.
En man och en kvinna på en skoter.
En grupp dansare med gröna skjortor håller alla hand i en cirkel, en dam har en vit skjorta.
Två kvinnor i svarta hattar står på gatan.
Solljuset kastar långa vertikala skuggor på baksidan av en unga flickors jeansjacka.
Tre kvinnor i blå och röda kläder bär en banderoll.
Fyra par som utför dansrutiner är färgglada gröna och vita kostymer.
En man lagar mat medan en annan vaktar.
En belagd medelålders man tittar genom ett teleskop på himlen på natten.
En man i en rutig skjorta tittar genom en teleskoplins.
Det finns flera personer på en båt och en är person som släpper sina lådor och mooking förbi.
En man i grön jacka som fiskar från toppen av en sten.
Polisen sätter gul tejp från en dörr till ett träd för att hindra åskådare från att komma in i området.
Mexikanska räddningsarbetare hjälper till att ta bort en man från ett kraschat fordon.
En brandman i uniform håller i en röd slang
Två män bär sin dotter på sina axlar.
En person med svart hatt och en facklig jackväska går på en trottoar passerade en gammal stenbyggnad, vars gröna fönster säger "mooch art".
Två personer som sitter utanför en glasbyggnad.
En man sitter på en bänk och pratar på en mobiltelefon medan andra går över en gångväg ovanför honom.
Invånarna ser efter efter en olycka mellan en röd och en svart bil.
Akutsjukvårdare, brandmän och poliser på platsen för en bilolycka.
En man använder en yxa för att göra gårdsarbete.
En grupp brandmän och tjänstemän förbereder sig för att svänga en bil höger sida efter en krasch.
En greyhound hoppar över gräsmarken.
En man i en svart och vit keps tittar in i en silverpontiac.
En trappa med gröna växter som växer på sidan.
Detta är en scen av en produktions besättning utanför på en gata nära en deli.
En brun hund har en lila skiva.
En man i orange röd skjorta tittar på två monitorer på ett skrivbord som också har sin fot och en Staples Easy-knapp på den.
Folk sitter i stolar längs en trädkantad trottoar.
Två kvinnor står på ett öppet fält, tillsammans med två hundar, en kvinna håller en hink, den andra en jacka.
Arbetare i hatt sveper löv nerför en gata.
Mannen bär svarta glasögon och v-neck t-shirt bär liten flicka i randiga byxor upp och ner.
En maskulin gentleman går nerför gatan och bär på en portfölj.
En kvinna bär en blå och vit randig skjorta medan hon sitter.
En man står bakom en jättegrön maskin.
En man sitter utanför i en blå gräsmatta stol och målar en man med svart hår på en duk.
Folk klättrar och vandrar nära en sjö.
En bil och många människor står på vägen.
Ett par kopplar av i en paddelbåt på en vattenförekomst.
En äldre kvinna i mörk rock håller ett paket papper hårt.
2 små flickor äter glass.
En ung kvinna i svart skjorta som går på en gata.
En man och en kvinna som håller ett barn går förbi några trämöbler.
Asianen i grön hatt och grön, orange och blå väst tittar på något.
En asiatisk kvinna i vitt förkläde och mask, med orange handskar tar en bild.
En man sitter på gatan under ett paraply med symaskinen och byter kläder.
Tre personer som bär vita hattar rider på en gaffeltruck.
En dam rider längs vägen på en motorcykel med en person med vit hjälm.
En man i svart kostym går.
En grupp på fyra barn går över gatan, när en vuxen tittar nerför gatan.
Två män med västar i kampsport.
En man, som bär en blå jacka, sparkar en annan man, bär en röd jacka.
Japanska människor som sitter i en riktigt tjusig café läsning.
En kvinna klädd i grått och en pojke klädd i en vit skjorta som leker med leksaker på marken.
En man i grön skjorta väntar medan polisen förhör några snowboardåkare.
Två män utövar kampsport en har sitt högra ben i den andra mannens ansikte.
En dam som håller en mikrofon stående på en scen.
En blond kvinna sjunger in i en mikrofon och ger "okej" symbolen med sin vänstra hand.
Man och kvinna håller räcke tittar bort i fjärran.
En arg man i en grön Seattle Seahawks hoodie lutar sig mot ett räcke.
Folk njuter av underhållningen på Summer Concert Series.
En man i hatt spelar en akustisk gitarr med ett band på en utomhusplats.
En kvinna målar ett tecken på en blå tegelvägg.
En ung man klädd i en blå jacka håller en staty över huvudet.
En man och en kvinna står på en scen.
En man med en rosa kamera som fotograferar en rockkonsert.
Ett band uppträder för Good Morning Americas Summer Concert Series.
En kvinna i en blå jacka läser en bok bredvid en annan kvinna som läser en tidskrift.
En man och kvinna som rider på en tunnelbanebil.
En man med en vagn går längs en vägg täckt av graffiti.
En vit hane spelar trummor.
Himlen lyser ett livfullt gult i solen.
En man i svart flyr med rep på balkongen.
En grupp människor möter mot en bro över vattnet.
Två unga kvinnor som messar med en cykel.
En folkmassa som blir vild när konserten tar slut.
En man balanserar en papperslykta på sin utsträckta hand.
Många människor står runt en gata bredvid en skylt
Man med Adidas gymväska går nerför trottoaren.
En äldre man som spelar ett instrument i regnet.
Ung flicka står i sin barnvagn på gräset.
En man med kamera och en annan man med barnvagn står i ett inhägnat område.
Tre kvinnor i svarta klänningar går nerför gatan
En överviktig person med sandaler läser en tidskrift på en bänk.
En man omgiven av tallrikar och tallrikar med mat.
Dessa tre flickor bär sommarklänningar och leker med hunden i gräset.
En man från Taiwan har ett tecken som protesterar mot regeringen.
En kvinna i jeans och en blå tanktopp som ligger i ett träd.
Två tjejer visar något för varandra.
En upptagen butik full av folk som handlar i butiken.
En kvinna med paraply sitter på en stenbänk.
En man hukar sig i gräset för att ta en bild av en blomma medan en smal kvinna tittar på.
En grupp musiker uppträder på gatan.
En skara människor står bredvid en nummer nio, antingen kliver på eller hoppar av.
En kvinna i en konstig uppsättning av kläder.
En man i militären går med sina två döttrar.
Två personer cyklar i stadstrafiken.
En ung svart pojke med randig skjorta, svarta shorts och svarta regnstövlar som ligger på en rad gula gatubarriärer.
En kvinna i vit utstyrsel går upp för trapporna.
En afroamerikansk man, lagar mat på vad som verkar vara en professionell matlagningsserie.
En äldre tungset man vilar på en bänk med sin kundvagn i närheten.
En man tittar på vad som verkar vara en kartong av en kvinna i ett kök.
En man med käpp går på trottoaren.
En grupp tonåringar sitter på trappan och tittar på en man och en kvinna.
Kvinnan går bakom två brevbärare droppar i gräset.
En afrikansk amerikansk arbetare som sätter mat i ugnen medan han tittar på kameran.
Ett barn som bär rosa sitter i en barnstol.
En man i röd skjorta och en blå hatt sitter på en trottoar och rör vid dricksglasögon.
En brunhårig kvinna lyssnar på en drink.
Två pojkar ler medan en kvinna ligger bakom dem i en barnvagn.
Två kvinnor bär mobiltelefoner och har ljusa klänningar.
En blå Harley motorcykel är en av en grupp motorcyklar som ägs av motorcyklister.
Kvinnan lagar skorna medan mannen tittar på sin mobil.
Två tjejer med vit dans på kvällen utanför.
Flickan i den grå skjortan har mycket mörkt hår.
En kvinna bär en grön tank topp och ovanliga halsband vid ett bord i en restaurang.
En kvinna i klänning och Capris lägger ut bilder
En dam i blå skjorta har en väska under vänster arm.
Kvinnan i lila skjorta stirrar i fjärran.
En man finner en unik plats att sitta och vila på en strandpromenad i staden.
En kvinna i vit skjorta går med en skjortlös, tatuerad man.
Dilapiderade byggnader i bakgrunden av en hel del grönt gräs.
Kvinnor som bär jeansjacka över randig skjorta går på dockgård
En kvinna med en mycket stor svart peruk och jättesolglasögon håller en spegel upp mot ansiktet.
En kvinna som står framför saker och ting.
En flicka sitter ner medan hon tittar på något.
En man tröstar sin vän längs gatan.
Folk går längs en strand med en brygga i bakgrunden.
En äldre man står ute på natten.
En medelålders man läser en plakett på ett träkors som ligger i ett fält med stängsel och träd.
En ung kvinnlig sprayfärgskonstnär arbetar på en målning.
En man som bär vit t-shirt och hörlurar använder sprayfärg medan han arbetar på en väggmålning.
Två tonåringar sitter på en brygga och kollar sina mobiler.
En grupp människor som cyklar och går över en väg i staden.
Folk väntar på att korsa en gata på natten.
Manlig surfare med gul surfbräda och hund går ner pittoresk strand och stora klippor.
Tre damer i kostym går genom ett köpcentrum.
En gammal man och kvinna på gräs mellan rader av amerikanska flaggor.
En kvinna håller en picketskylt på en trottoar.
Kvinnan kollar apparaten när hon trampar ner på gatan.
Ett stängsel skiljer en kvinna som håller en röd flagga från en polis.
En man som går genom en livlig stad där en annan man på en cykel transporterar varor.
En kvinna och två barn förbereder en drake.
Tre kvinnor är ute och dricker tillsammans.
Asiater som står i ett företag.
Lycklig ansikte av människan talar i mikrofon som hålls i handen framför tegel byggnad.
En äldre konstnärsmålning medan hans sittande hund tittar på.
En man i svart och vit rutig skjorta sitter vid ett bord i restaurangen och beställer mat.
En man i vit skjorta som tar en bild.
Två kvinnor går mot en brandpost, målad med ett ansikte på.
En svart kvinna som håller i ett paraply korsar gatan.
En grupp kvinnor i sportuniform spelar frisbee på ett fält medan andra tittar.
En gatuartist målad i guld står av en guldtäckt gammal tidskamera.
En baseballspelare försöker märka ut en löpare.
En kvinna fifflar med sin telefon på ett matställe.
En kvinna går nerför gatan på sin mobiltelefon medan hon håller en kopp kaffe.
Tre män står bredvid varandra och bär olika färgade skjortor.
En man med röda glasögon och lockigt hår står på en livlig gata.
En man går på en smal gångväg.
En man i en grå tröja som gör ett ansikte medan han spelar trummor.
En person som bär rullskridskor åker skridskor längs ett räcke.
En man i rullskridskor sitter ner på en utomhusåkning park.
Tre personer går förbi en väggmålning av en ko.
En grupp människor samlades i ett stort rum med vackra arkitektoniska element.
En mor och hennes två döttrar stannar på en gårdsplan.
Den blinda kvinnan i den rosa skjortan pratar med en man utanför caféet.
Kvinnan på gatan håller en Starbucks kaffe.
En man som bär sina traditionella etniska kläder skrattar när han ser en show.
Folk går runt elefantmodeller för bebisar.
En motorcykel racer i en blå och rosa kostym gör sig redo att tävla.
En man i paraplyhatt sitter nära ett palmträd bakom en grupp shoppare.
En man sitter ner klädd i blå handskar och bär en vit jacka.
En kvinna går en hund i koppel.
En person som ligger utanför och läser en bok under dagen.
En kvinna springer i ett lopp medan åskådare hejar på henne
Mannen sitter på röda trappsteg utanför lägenheten med röda dörrar.
Två personer går bredvid en vägg med graffiti.
En smal man och en stout man går på en strandpromenad.
En hona som ligger på magen i vattnet utanför med paraplyer.
Två unga damer sitter på trappan till en rustik byggnad.
En man står bredvid en polisbil.
En ung man som bär grå skjorta står utanför ett timmerhus medan han ler.
Folk sitter vid ett bord medan en man pratar med en mikrofon.
En stadskorsning med en man på cykel och en butik på hörnet kallas SWATCH.
En livlig gata med shoppare som tar sig hem.
En man i grå skjorta står utanför tunnelbanan.
En baseballspelare ger sig ut på en boll.
En man i blå skjorta som sitter på en blå stol.
En kvinna i jeans som går med ett paraply.
En man i röd skjorta och vita shorts går bakom en man i vit skjorta.
Flera asiatiska människor är på ett tåg.
Flera personer sitter på platser nära ett litet bord med drinkar.
En kvinna tittar ner från en hög punkt ovanför ett lugnt blått hav.
En brun hund hoppar över en kedja.
Två män sitter på en trappa bredvid nummer fem.
Medan en man med grå t-shirt dricker en koupé av röda stripe öl, talar en man med en grå t-shirt till en annan man som bär en blå knapp upp skjorta.
Kvinnan bär en blomtryckt skjorta.
Detta fotografi fångade en man och en kvinna som åkte skridskor i en sammanflätad pose.
En grupp äldre män och kvinnor sitter och lyssnar uppmärksamt i fällstolar av metall.
Det finns en stor skara människor med paraplyer.
Fyra män i gröna uniformer sopar upp gatan efter en parad.
Två män spelar didgeridoos framför en eldstad medan en sibirisk Husky ligger på en soffa.
Man på sopbilen jobbar hårt för dagen.
En kvinna står framför en vägg med en massa graffiti.
En leende konstnär knäböjer på trottoaren.
En man i en ljusblå skjorta är böjd över att justera sin känga, medan hans hatt ligger åt höger.
En grupp människor i en återförening diskuterar ett mycket viktigt ämne.
En man i khakis och en blå skjorta talar in i en mikrofon inför en grupp.
Man och kvinna pratar på seminariet.
En medelålders man som bär en blå huva och en rutig hatt står med uppvikta armar utanför en stadsbyggnad.
En grå "labradodle" hoppar över en annan stor hund.
Tre män sitter, och en man står, på baksidan av ett fordon.
Mannen i de röda shortsen har en tatuering på benet.
Två barn står mot en tegelvägg i solljuset.
Hon går förbi den vackra blå väggmålningen.
En man i glas med öl och eld
En arabisk kvinna blir intervjuad av pressen.
Gul taxihytt som rör sig över bron och stora byggnader i bakgrunden.
En gammal man spelar gitarr.
Två unga kvinnor håller händerna nära ett träd.
En skyltdocka klädd i underkläder annonseras.
En man lägger sand på marken nära en stor stadga för en dam som sitter ner i en röd klänning som håller en flaska.
Folk äter på en restaurang.
Detta är ett fyrvägs stopp med tre bilar, en cyklist och två fotgängare.
Det är en man som går på trottoaren.
Två män, den ene klädd i röd skjorta och svarta byxor och den andre klädd i vitt, spelar basket utanför en tegelbyggnad.
En brandman som står ovanpå en brandbil.
En häst har störtat i en arena och ryttaren kommer ut från ryggen mitt i luften framför en folkmassa i läktaren.
Många människor går upp och ner ChinaTown, möjligen under en händelse.
En ung pojke som bär en svart och röd klänningsskjorta ryser när han tittar bort.
En man som säljer en bunt ballonger på en strandpromenad
En stor grupp människor stiger upp i en trappa och lämnar ett rum med orientalisk skrift i taket.
Folk har någon slags dag rättvis.
En man i en blå randig skjorta och jeans tillsammans med en kvinna i en brun skjorta som går tvärs över gatan.
En tungsint man med två rödhåriga bebisar i knät.
En grupp människor står bredvid en "ingen lastbil" skylt och en gul gatuskylt.
En mörkhyad liten pojke med hörlurar i.
Fyra personer är på en röd bro med ett rör som går över den, en del går medan en del står på plats.
En kvinna med rakt blont hår pratar på en mobiltelefon utanför.
En offentlig samling av olika slag som huvudsakligen består av människor av afrikansk härkomst.
Fyra män står utanför nära en vit lastbilssäng.
En grupp tjejer runt ett bord fullt av tyg.
1950-talets polisbilar på matbilen.
En blond dam i en dekorerad blå klänning täcker sitt ansikte med handen.
En man använder en hammare och mejsel för att göra skulpturer.
Gatan i Europa där en grupp män sitter på sina motorcyklar.
Två män i en gul Penske lastbil
En person i svart lutar sig mot en byggnad i en strimma av solsken.
Skäggig man i stringtrosor pratar med kvinna en solig dag.
Cityscape med fyra män på cyklar som fungerar som fokus för bilden.
Ett gammalt par som gick nerför en gränd och höll varandra i handen.
Unga damer som jobbar på sina datorer, studerar och kopplar av samtidigt.
Två män förbereder sitt dryckesstånd.
En blond kvinna i en blå tank topp tittar på en oidentifierad figur framför kameran.
Tre kvinnor passerar förbi en affisch på gatan.
En kille i shorts och en baklänges mössa målar en vägg utanför.
Två personer, en sittande och en stående, framför en graffitimålning.
Två boxare landar samtidigt på varandra.
En man drar en skottkärra lastad med tegelstenar.
En kvinna i svart hatt och svart skjorta som står framför en Red Bull Car.
En brunett dam i en blå skjorta ringer upp en kund i en butik.
En cyklist med grön ryggsäck och hjälm på gatorna.
En grupp människor tittar över avsatsen.
En man klär sig i en militäruniform tittar genom ett mikroskop medan en skallig man i vit rock ser på.
Tre små barn i ett öppet fält tittar mot himlen.
Kvinnan i svart klänning med blommor tar en bild på konstmuseet.
En man i brun kostym går nerför trottoaren.
En kvinna i grön skjorta som svingar, med bara en sko på.
En lärare som undervisar sina elever i klassen.
Två kvinnliga arbetare i hattar som serverar mat från ett stall.
Den här personen klättrar upp på sidan av ett berg.
Männen i den långa klädgarderoben håller på med en show.
En klättrare som stiger uppför ett berg
En kvinna i blå skjorta målar två fönster med gröna nyanser.
En man i hatt som ligger ner medan han fotograferar.
Personen lägger sig på en orange duk framför en jättestor affischtavla med gating framför den.
En man i grön skjorta står bredvid en bil på gatan.
En man som står framför en pizzarestaurang med lådor framför.
En man i en färgglad slipsfärgad skjorta går förbi en nagelsalong.
En grupp professionellt klädda människor sitter nära varandra är ett centrum av en stad.
Människor samlas utomhus på natten.
En man i en ljusgul skjorta som står utanför en ljusgul byggnad nära en telefonautomat som har en ljusgul handset.
En afrikansk amerikansk man står framför en brandstation i Harlem.
En man i vit skjorta står framför en klädaffär.
Bicyklisten tittar åt höger när han färdas genom trafiken.
Kvinna i blå klänning och bär en svart handväska, rider en scooter nerför gatan.
En äldre man i en rutig skjorta som lutar sig mot en restaurang.
Byggarbetare tittar på från toppen av byggnaden medan ytterligare två är upphängda från en kran i en korg.
En kvinna dricker en öl medan hon tittar på en utomhuskonsert.
En grupp människor med färgglada flaggor i centrum.
Folk i svarta hattar samlades i centrum.
En ung kvinna hoppar upp i luften med USA:s Capitol byggnad i bakgrunden.
Folk rider motoriserade vertikala skotrar längre ner på gatan.
Folk som sitter på marken och ser på när en liten pojke och en man gör något.
Flera människor rör sig bort från ett färgstarkt torn.
Tre unga män tittar på en tennismatch på en stor skärm utomhus.
En man är ute och hackar mat på ett bord.
En man i röd skjorta som håller en käpp beställer lite mat på marknaden.
En kvinna som håller i en dryck går nerför gatan.
En man med vit skjorta och tatuering sitter inne i ett glassställ täckt med bilder av läckra godsaker.
En man läser en bok, på en trottoar, medan en kvinna väntar och andra fotgängare går förbi.
En polisman pratar med flera män på en livlig stadsgata.
En kvinna i rosa klänning sitter på en cykel.
En kvinna i en blå skjorta som sitter vid ett bord med sin anteckningsbok, penna och laptop.
F.d. guvernör i New Mexico, Bill Richardson i Mellanöstern håller tal.
En man i vit hatt, solglasögon och mörk skjorta talar in i en mikrofon.
Stor man i svart skjorta bredvid polis som går iväg från mannen i blå skjorta och ryggsäck
En kvinna står i en vit lastbil och sjunger medan folk tittar på henne.
En grupp människor protesterar i en stad.
En kvinna med huvudbonad och traditionella kläder läser in i en mikrofon från ett papper.
En grupp låter sin politiska åsikt bli känd.
En liten pojke som bär hjälm ler medan hans far gör lite justeringar på ryggen.
En man i svart skjorta som lastar eller lossar en blå honda.
En grupp människor väntar på trottoaren, klädda i hattar.
En grupp av Mellanösterns arv marscherar nerför en stad gata protesterar.
Det är många människor som deltar i en parad liknande aktivitet på gatan.
En man i en restaurang som man tittar på genom ett fönster.
Flera män och kvinnor protesterar mot Israel medan en man i en blå skjorta skriker åt dem.
En skara människor marscherar.
Ett band som spelar en konsert framför en måttligt stor publik
Tre människor sitter och väntar.
Två män står på trottoaren med sina instrument på ryggen.
En fotograf fotograferar en utsmyckad byggnad.
Två kvinnor och en man står framför en målning av Cher.
Folk står i kö vid en lastbil och väntar på att få köpa glass.
Två personer rusar över gatan medan regnet faller från ovan.
En grupp människor sitter på en stenig strand.
En polis med en kirurgisk mask på står framför en grupp flickor i uniform.
Folk går nerför en gata i ett obefolkat område.
En motorcyklist stannar vid en tom crosswalk, medan trettio eller fyrtio motorcyklar och cyklar sitter parkerade på gatan bredvid honom.
Tre arbetare är ute på natten och jobbar.
En man i vit skjorta läser en tidning.
Ett par njuter av landskapet medan en fotograf fångar det på film.
En molnig dag i en stad håller inte folkmassor av män och kvinnor borta på trottoarerna.
En asiatisk flicka modellerar gummistövlar.
En man med röd keps och tröja står bredvid en äldre bil och stirrar på en ung, blond kvinna när hon går förbi.
En affärsman i soldräkt sover på trottoaren nära en byggnad.
En liten flicka som rider en tvåhjuling, bär sin hjälm nära gatan med förbipasserande bilar.
Två kvinnor med svarta t-shirts sitter i gräset.
En tjej med blont hår med en ärmlös topp hålls fången av en kvinna.
Mannen går lilla flicka med ryggsäck tvärs över gatan.
En kvinna med rött hår går nerför en trädkantad stig med en brindled hund som följer henne.
En tjej i vit jacka säljer bakverk ur en låda.
En man i en babyblå arbetströja pratar i telefon på den livliga trottoaren.
En kvinna i en blå tank topp och blå byxor joggar.
Tatuerade kvinnliga hipster med överdimensionerade bälte leenden medan en annan kvinna står i bakgrunden.
En man med glasögon bär en skjorta som säger att man ska åka till centrum.
Två svarta män i svarta rockar går längs gatan med kvinnor som tittar på dem.
En skara människor i ett utomhusområde.
En man i vattendräkt med ett äpple i handen tittar över en klippa.
Två personer sitter i hattar och nyanser.
En man med brunt hår som spelar trummor.
En kvinna på en ljus gata spelar fiol.
Ett par går genom ett hektiskt område med många människor.
Folk som står på en station.
En kvinna i svart skjorta och shorts går genom en fontän.
En man som röker och håller kopplet mot en hund står bredvid en kvinna som bär solglasögon.
En tjej i blå klänning och en kille i jeans går in i en butiksfront tillsammans.
Kvinna med långt hår på cykel tittar på ett barn.
En liten flicka, vid ett staket, ser ut som hon pratar på en mobiltelefon.
En man som bär rutig hatt sitter i en fåtölj och läser en tidning
En kvinna med mörka kläder och en hästsvans som går förbi ett metallstängsel nära en busstation.
En ung kvinna går ensam genom en bussterminal.
En kvinna i röd klänning står bredvid ett stort träd.
En äldre herre förbereder sig för att träffa en golfboll.
En man med mörkblå skjorta och hatt bär glasögon bredvid en taxi.
En man som bär en röd rutig kilt som står framför ett förbipasserande barn.
En kvinna i röd kjol med blommor går nerför gatan.
En ung pojke i hatt fiskar ensam.
En silverbil som kör förbi ett hotell där folk står utanför.
Två damer skrattar på gatan.
Vissa människor sitter på en järnväg över en sjö.
En ung kvinna som går på en livlig gata
En tjej med uniform stående på trottoaren med något rött och blått i handen.
De här två kvinnorna är på Giorgio's och har kul.
Två hundar med huvudet nerför ett hål och deras svansar sticker rakt upp.
En liten asiatisk pojke som äter pizza.
En asiatisk kvinna håller i ett stort blått och vitt rör medan hon tittar på en annan kvinna och en röd buss passerar henne.
Man bär svart skjorta kastar en yxa.
En fullsatt gata, i ett asiatiskt land, där byggnaderna domineras av Seiko-byggnaden.
De unga pojkarna vid bordet spelar ett spel.
Två små barn sover på en soffa.
En scenkonstgrupp deltar i en liten parad.
En pojke som leker med bollen i huvudstaden Berlin, Tyskland, i Europa.
Två män med ryggsäckar på att titta på underkläder i ett fönster.
En äldre kvinna lutar sig mot balkongräcket i ett hyreshus; hon tittar ut över en gatulampa.
En hund springer längs havets surfing.
En kvinna i underkläder på en kudde medan män tittar på henne.
Två fashionabla tjejer står på en trottoar framför vissa cyklar.
En ung pojke i en röd flytväst simmar i en pool.
Två unga flickor går i en parad.
En tunnelbanescen, med ett blått tåg som rör sig genom stationen medan passagerarna går och väntar runt.
Korstågen marscherar längs vägen.
En man med beigeskjorta har hukat sig ner på gatan bredvid några huggna stenar.
En bil med stora väskor på toppen.
En kvinna springer framför en randig vägg.
En man rider en jetski över havet.
Ett par i en stad där turister besöker, men de är olyckliga.
En man sprintar av en annan man med ett paraply.
En man målar en annans ansikte vid ett utomhusevenemang.
Ett par kyssar utomhus, medan ytterligare ett par tittar på.
En man i svart skjorta och jeans går vid havet.
Den urbana trolly's av en stad på en solig dag.
En man i panamamössa och flygarglasögon samtalar med en annan man i en grå sportrock och jeans.
En gatuvy med bilar och byggnader.
Ung blond flicka ser osäker ut när hon matar färgglada fåglar utanför.
En liten flicka som ler i en färgglad stickad hatt.
En man som fotograferar en bro på floden under solnedgången.
En grupp räddningsarbetare övervakar en kraftig försämring på en gata i staden.
Folk samlas utanför en byggnad där 'Love Story' hålls.
En kvinna och ett barn som gör en varelse av pappersprodukter.
En man i vit skjorta och en kvinna i röd skjorta dansar utomhus med många människor runt omkring.
En grupp människor tittar på varor på ett bord.
Flicka i färgstark topp och höga klackar dans
En man i en blå skjorta som målar något utanför.
En vuxen man håller i ett manligt barn som tittar på ett djur och en vuxen kvinna håller ett kvinnligt barn.
En svart och vit hund springer genom ett kofält.
Framsidan av en matförsäljare i en park.
En kvinna som målar något på en liten flickas ansikte.
En man i röd rostfärgad rock som bär en stor träpåle.
Grupp av asiska män som spelar volleyboll
En kvinna i orange skor som röker och läser på en parkbänk.
En gammal asiatisk man som stod i dörren till en byggnad.
En man i khakijacka och keps går nerför gatan.
En man i blå skjorta går nerför en trottoar.
En man som bär hatt går och bär en stolpe med en krok i ena handen och en stor aluminiumburk i den andra.
Carnival Barker står framför ett cirkustält.
Härlig stadsscen som visar en klarblå himmel, tre gamla byggnader och en smal gata med järnvägsspår.
Fem soldater håller och siktar sina vapen.
En soldat skjuter när han står bredvid en vägg.
En grupp människor med utsikt över vattnet från en båt.
Det finns en individ i denna bild med en hård hatt om och en radio i handen verkar vänta på instruktioner.
En soldat hukar sig bredvid sitt pansarfordon parkerat under en bro.
Fyra personer i nöddräkter och hjälmar sprutar vatten bakom en cementvägg.
En soldat som duckar och håller i ett vapen med gröna kläder.
Två brandmän släcker en brand vid en soptipp.
En militär man kikar ut från toppen av sin stridsvagn.
Den unge mannen med en vit tröja går bort från den vita Acura bilen.
Två män går tillsammans längs en trottoar.
En man och en kvinna undersöker färskvarornas varor i en livsmedelsaffär.
Kvinnan i rosa skjorta och svart kjol går nerför gatan.
En gammal man knuffar en vagn förbi en skoaffär.
En man som går längs gatan och bär på en sopsäck.
Två flickor går nerför en asfalterad trottoar i en stadsmiljö.
En liten bebis som bär blå kläder tar lite frukt.
En grupp soldater står med vapen framför ett pansarfordon.
Tre män i militäruniform håller i vapen.
Två unga militärer i kamouflage med automatvapen.
Polisen ser ner på ett gevär i Thailand.
En ung kvinna som stod på däck på en båt och stirrade på sin mobil medan hon satt på vattnet.
En kvinna med blommössa sitter bakom en man vid piren.
Brandmännen på bilden gör sig redo att använda sin brandutrustning.
Brandmän sprutar in en slang i en brand.
4 Brandmän som använder en brandslang för att släcka en brand.
Beväpnade styrkor går i ett område fyllt med skräp.
Brandmän satte vatten på en rykande hög med skräp.
Två soldater tar sin tillflykt bakom några skyddsräcken.
En grupp armémän och kvinnor håller vapen och springer nerför gatan.
Kvinna med paraply ridning cykel bakom par promenader medan du använder ett paraply
En gammal dam står bredvid en antik i en klänning.
En man som jobbar på en vävstolsliknande apparat.
En man som bär vitt hänger tråd på en stolpe av bambu.
Fyra kvinnor med tatueringar håller små flaggor.
En stor grupp människor samlas på en innergård, med en del som ligger på mattor.
En vit hane pratar på en mikrofon.
En hund biter ett föremål som erbjuds av en person.
En grupp människor står utanför.
Många vita står bakom flaggor och en banner, bredvid stora grå byggnader.
En person spinner bomull i tyg.
Folk går på en stadsgata och en man som håller en gul flagga.
En grupp på fyra personer sitter på en stenmur.
En grupp barn som står på en scen och håller gula klockor och pekar på något.
Två arbetare möter varandra i gröna kläder.
En grupp på 70 eller 80 år kaukasiska män och kvinnor satt och hade en diskussion.
Stor publik på en Birmingham händelse.
En clown med gul peruk och skjorta och flerfärgade hängslen håller en orange ballong i båda händerna medan ett barn i svart hatt ser på.
En massa människor, med en man som kollar sin telefon mot dig.
En man som har två broschyrer poserar på en upptagen NY-gata.
Två kvinnor njuter av de öppna landskapen i en park.
Folk går i en parad, som andra tittar på.
Föreställare i färgglada kläder står på en scen.
En ung pojke med röd ryggsäck och blå skjorta har utsikt över landskapet av ett historiskt landmärke.
Två kvinnor håller en röd och vit flagga medan två andra kvinnor tittar på.
En stor grupp i rött vitt och svart uppträder på en scen.
En grupp människor uppträder tillsammans på scenen.
En skara människor håller vita flaggor med röda kors.
En man står och håller tal på en scen.
En kvinna i en blå och grön klänning står framför en kvinna i en lila klänning med en vit spetskrage.
Människor, några i uniform, mala omkring på en gata.
Två asiatiska kvinnor står bredvid ett bord som har mat på sig.
En stor grupp människor tävlar genom en kraftigt trädbevuxen park.
Ett maraton börjar på en stad gata under en JP Morgan banner.
En polis bevakar ett maraton.
En man är ute med sina små söner, och kysser en medan den andra leker.
En grupp campare vid sjön, tillreder och grillar mat
En svagt klädd ung kvinna driver en mountainbike på en rekreationsstig längs en vattenförekomst.
En ung person skateboards av den färgglada väggmålning målade på byggnaden.
En man i vit skjorta spelar saxofon på en scen.
Hundratals människor springer ett maraton genom en stad.
Många vakter står framför startlinjen för ett lopp.
En massiv krona väntar mitt i staden.
En grupp människor står runt en lång rad bananer.
En man som går längs sidan och städar upp.
En maskerad läkare som bär glasögon utför en operation.
Stor ljusfixtur i fullsatt operationsrum.
Läkarna försöker genast reparera den läckande hjärtklaffen.
En man sitter i ett vitt rum bland olika vetenskapliga maskineri.
Fyra män och en kvinna sitter bakom ett bord, medan ett hjul sitter på väggen i bakgrunden.
Tre män klädda i operationskläder opererar en patient.
En kirurgisk RN i blått skrubbar kontrollera inställningarna på maskinerna före operation.
Två kvinnor som bär cowboyhattar går nerför en trottoar och bär påsar.
En man i hatt sitter vid ett av flera bord inne i ett skärmat tält och tittar på människor som går förbi utanför.
Tre personer går på en strand.
En man med svart skjorta och mikrofon utför en demonstration vid ett evenemang.
Två små hundar sitter nära ett träd.
En flintskallig man får sina skor tvättade i ett gathörn.
Ett par sitter i parken nära ett litet vattenfall.
En del människor går uppför en trappa nära vattnet.
Tre kirurger som opererar en patient.
Ett läkarrum med en man klädd i blått.
En person är i ett operationsrum.
Två män i kirurgklänning slutför en operation i en operation.
Ett operationsrum fullt av läkare och sjuksköterskor.
En grupp kirurger som bär skrubb utför en operation.
En kvinna håller ett barn i gräset
Medicinsk personal ser på som en medicinsk procedur sker på en videomonitor.
Läkaren observerar en bild före operationen.
En grupp läkare som utför en operation i en operation.
Läkare med skyddskläder opererar.
En man som väntar på läkarens order att operera en cancerpatient på operationsavdelningen.
Några turister besöker ett landmärke.
Den bruna och vita hunden bär en käpp i munnen.
En kvinna i en vit blus står framför en skara sittande barn.
Musik kan skapas, genom blåsinstrument, med blåsinstrument, och de är alla avnjutna av olika folk, över hela världen.
Tittar på en gata med en skylt ovanför butiker som säger Välkommen till Golden.
Två män hoppar i luften för en bild.
En hund som simmar med en käpp i munnen.
Indiska kvinnor i färgglada Saris tala och titta igenom material medan ett barn sitter i närheten.
En man med hatt vänder sig om och tittar på kort.
En liten pojke bär en t-shirt som säger att Gidday tittar upp mot himlen medan han njuter av ett mellanmål.
En naken cowboy som fotograferar med två damer.
En uppsättning nycklar i låset på en öppen låda på en utvändig stolpe.
En flicka tittar ner i en pool under en fontän.
Två hundar med rosa hår har koppel.
En man med orange ryggsäck i ett buskigt område.
Det finns många människor på den här livliga asiatiska gatan.
En livlig gata har flera människor runt omkring och cyklar radas upp i rad.
Några få människor står utanför affärerna i en asiatisk stad.
En samling unga kvinnor på en orientalisk marknad.
Två män, en med flera tatueringar på axeln och överarmen, går på en trottoar täckt av tuggummi.
En man i idrottskläder som håller en vattenflaska i gång.
En vandrare står på en kulle och tittar i fjärran.
I Italien är gatorna fulla av människor.
En man och kvinna går på en restaurang som har skyltar på kinesiska.
Två kvinnor låg på magen i solen.
En man i skinnrock väntar med en annan vid en busshållplats.
Två asiatiska kvinnor sitter i skuggan under ett träd.
Fotgängare som går på en fullsatt gata i en asiatisk stad, sett från baksidan.
En grupp människor väntar på en tågstation.
En äldre man sitter bredvid sina skor och jacka medan han lutar sig mot en vägg.
Ett leende ungt par promenerar arm i arm nerför en Paris gata.
En kille med långt hår och stor mage som går vilt förbi en väggmålning av en tjej som ser galen ut.
En publik är runt en showgirl som bär en vit huvudbonad.
Två hundar är lite ovänliga med sina ägare som sitter ner framför en tid realty tecken.
Folk tittar ner på något bredvid en stor stenbyggnad.
En man i blå skjorta funderar på vilken bok han vill köpa.
Unge man som sitter vid en fontän i telefonen.
Många människor i röda sporttröjor går och pratar på en stad gata.
Ett par människor går nerför en gata upplyst av skyltar på natten.
Det finns en ung man på en skateboard framför ett matbås.
En kvinna med barnvagn går mot en grupp unga män.
Tre barn leker med en gul leksak på en grön kudde.
Många cyklister och andra människor på en gata
En grupp av tre unga flickor i klänningar går längs en gata.
En man i en rutig skjorta blåser i ett horn.
En kvinna som håller en liten flicka i handen och går över en bro.
En man läser tidningen medan han dricker.
Två unga pojkar som använder sparkbrädor för att lära sig simma.
Barn som leker i en pool med rent vatten.
En gammal man med kostym, slips och kaptenshatt står mitt ibland folk, med en arg blick i ansiktet.
En kvinna står på trottoaren, framför en korsning.
En man i svart klänning går nära en affisch på en plattform.
Vissa människor nära en vattenförekomst med ljus överallt.
En äldre man med en vandrare som går framför en färgglad vägg, med flera saker på gång.
En flicka med mobiltelefon står under en gatuskylt.
En liten pojke med blå vantar som går över en trästigsbro.
En kvinna och en man som spelar gitarr medan en brunhårig kvinna pratar i telefon.
En person i ett rum inspekterar någon form av utrustning.
Flera kvinnor med långt hår och mini-klänningar går tillsammans.
En man står i dörröppningen medan en annan man går i ett rum som är i dålig form.
Damen i de vita byxorna har handen mot munnen.
En man i en blå mössa med en blå tröja pratar på en mikrofon medan en man utan skjorta ler.
En man arbetar på en grönsaksmarknad, med priser som visas i närheten.
Det finns många familjer som säljer olika varor, inklusive kläder, i en park.
Ett par som bär kimonor går längs en skuggig bana i Japan.
En man med röd väst som tittar på en man med orange skjorta som håller i en spegel.
Två man lutar sig mot en tegelvägg utanför
En äldre svart man spelar elgitarr på en gata.
En man i blå jacka står på en marknad.
En kvinna klädd i vitt och klackar går framför en vägg med en väggmålning på.
Smickrande kvinnor i en lila skjorta som kör ett lopp.
Två personer klättrar steg som leder till tre sammankopplade gröna statyer.
En man visar upp sin utrustning för åskådare.
Kvinnorna tittar på de vackra smyckena.
Två kvinnor kedjade ihop, en i röd klänning, den andra i blå skjorta.
Det finns en person som kör en lång cykel, framför en lila buss.
En kvinna i vit t-shirt, vita shorts och solglasögon.
En trång orientalisk marknadsplats på en smal gata.
En moderiktig ung kvinna som går genom gröna hus.
En man i en minikjol som försöker springa genom ett fält.
En kroppsbyggare som bär en Nike-skjorta kastar ett tungt föremål.
En man som bär kilt står på ett fält omgivet av flaggor och blommor.
En man och en kvinna står tillsammans vända mot varandra.
En man i jeansjacka målar ett tecken.
En man och en pojke tittar på vykort.
En skara människor på en gata nedanför en målad glasskylt.
Natten vid flodkanalen är upptagen.
En dam klädd i en vit, kort klänning bredvid ett bord dukat för två med en stenpir i bakgrunden.
En ung pojke som bär väst sitter omgiven av och leker med Legos.
Leende män som bär siffror som fästs vid deras bröst ras går nerför en våt gata.
Fotografer tar bilder på en flicka som sitter på en gata.
Det finns en åkare som bär en gul topp på sina knän på rätt spår.
En grupp kvinnor deltar i en roller derby spel.
En byggarbetare i overall och en gul bygghatt skyfflar smuts till en skottkärra.
En ung man tilltuggar medan han på en brygga tittar ut i en vattenförekomst.
En asiatisk flicka i en keps håller i en vattenflaska.
En man i röd skjorta och blå hatt fiske.
Flera människor tittar på andra spela inne i en uppblåsbar mån studsa karneval attraktion.
En pojke i randig skjorta som håller upp en fisk på en lina.
En skjortlös man som sitter på en bänk fioler med något i handen.
Turisten tar bilder på den vackra platsen.
En tjej med svarta byxor är att sänka en kamera på löpbanan.
De här kvinnorna åker skridskor i Roller Derby.
Tre kvinnor i matchande svarta och gula klänningar och en kvinna med orange hår.
En man med en stor kamera fotograferar.
En grupp tjejer som spelar roller derby medan en publik tittar på i bakgrunden.
Två män sätter upp ett hopphus.
En pojke i gul skjorta rider på baksidan av en annan pojkes cykel nerför en asfalterad gata.
Ungar fiskar i en sjö med sina fäder.
En man som bär förkläde ser en pojke arbeta på en cykel, och de är omgivna av andra cyklar.
En ung flicka fiskar i en sjö.
En man med skägg och röd hatt sätter sig ner med en drink i en papperspåse.
En matvagn körs nära en uteservering.
Tre kvinnor klädda i svarta kjolar och bh-toppar verkar ha börjat eller avslutat en dansrutin.
En gammal cadillac och en vit motorcykel på en gata.
En pojke cyklar förbi en grind med metallkyckling på.
Två kvinnor röker när de går på gatorna.
En grupp soldater marscherar i en parad.
En afroamerikansk kvinna som tittar på en affisch.
Den här kvinnan verkar gå på sidan av ett ljusblått hus.
En kille som tittar på stadskartan.
En äldre gentleman och en dam tittar på något som inte syns på fotografiet.
Två vuxna leder ett dussin barn längs trottoaren.
En liten flicka bär en rosa skjorta plocka upp små svarta objekt med en vit spade.
Tre kvinnor pratar och ser sig omkring.
En flicka i grön skjorta poserar humoristiskt med en cykel på en parkeringsplats.
En kvinna sitter på en sten vid vattnet.
En man sitter i en stol vid poolen och spelar gitarr.
En tjej med blont hår och en svart jacka som går längs en trottoar.
En kvinna nafsar på ett matföremål i sina händer.
En mamma och hennes dotter sitter i stolar på trottoaren.
En man hänger från en vågrät stolpe, som sitter i en byggnad, med en hand.
Kvinnor tävlar i en omgång roller derby.
På en smal gata kantad av hus, några med röda markiser, talar en man på sin mobiltelefon.
En kvinna och en man som sitter på en bänk framför en restaurang.
En man i vit skjorta läser ett papper medan andra sitter på en bänk.
En skara asiater som går runt i staden.
Tre kvinnor, med långt, okammat hår, står tillsammans, framför en stenvägg med peep-hål.
Folk står i ett gathörn i Asian City.
En man klädd i glasögon och en spetsig gasmask blickar i ångest och ilska.
Fyra tjejer i en pool som gör sig redo att hoppa i.
Ett stort antal människor samlas runt en vattensamling.
Två kvinnor står framför en karta.
Mannen sitter på bänken med en resväska framför skylten PADDINGTON.
En kvinna som står på en lutning med en röd väska.
Tre personer sitter tillsammans och konsulterar en anteckningsbok medan en man står och vakar över sina axlar.
Två män på hästryggen som en annan man kastas från sin böljande häst.
Unga flicka i en ljus rosa skjorta justerar sin kogirl hatt
En man som pratar på sin mobil på gatan.
En man ler ner från toppen av en totempåle en solig dag.
Ett litet barn som sitter på en bänk och äter något rött.
En kvinna med lila topp dricker direkt från en svart flaska.
En grupp människor som stänker i vatten.
Två män i hulakjolar står på toppen av en ramp i en lastbil.
Fyra män på kaffe, te och varm choklad.
En kvinna med en ljus orange ryggsäck står framför en trappa.
Damen pekar på sina kläder i torktumlaren.
En man i ett vitt förkläde håller en kyckling ovanför en stor gryta eller hink.
Två pojkar sitter och läser serietidningar.
En man med glasögon som står på en stege och målar en vägg.
En man som ligger på gatan.
En man i svart och blå jacka spelar en spelmaskin.
En kvinna i en brun puffig jacka går över en livlig gata.
En kvinna tittar på en röd halsduk från en av försäljarna på gatan.
Fyra damer tar en promenad.
En svart kvinna klädd i tanktopp och jeans håller ett koppel till en brun hund.
En kvinna med långt rosa hår sitter på en betongplatta.
Unga män springer på stranden för att träna för fotboll.
Folk står och tittar ut genom fönstret för att se berget.
En svart kvinna i gul och grön klänning som går längs en väg och bär en buske med en stor säck på huvudet.
Två flickor rider nerför gatan på enhjulingar.
En kvinna med en lång svart hästsvans och en flytande vit klänning.
En kvinna i lila topp bär ett rött och vitt paraply.
En man med en kamera runt halsen kör en moped i ett latinamerikanskt land.
En flintskallig man som står med handen i byxorna.
En äldre man i en rutig skjorta och jeans tömmer en kaffekopp i en soptunna.
Ett barn som bär en randig tröja trycker på en leksaksvagn.
Den lilla leende pojken lyfter pappret från presentlådan för att se vad som finns inuti.
Sju män klädda i orange skyddshattar arbetar på järnvägsspår.
Folk går i en byggnad där mat säljs.
En kille som sitter i en stol på gatan bredvid sin hund.
Två män i ett konstbås pratar med varandra.
På en öppen marknad inspekterar en man några vattenmeloner till salu.
Den här mannen ligger på trottoaren under graffiti på en vägg.
En hemlös man läser en tidning.
En man klädd i svart skjorta med djävulsögon som håller i två stora köttbitar.
Fem barn med hattar leker i leran på stranden.
Två barn står på en strand och gör ansikten, deras underarmar täckta av lera sträcker sig mot betraktaren.
En talare i ett klassrum.
Tre kvinnor ber med händerna vikta.
Två blonda kvinnor kramar varandra.
En grupp människor utanför en restaurang i ett inomhus shoppingområde.
Kunderna går omkring i en mataffär.
Två skateboardåkare går nerför en trottoar framför många parkeringsskyltar.
Två män håller skateboard och en man skateboard.
En ung man dränks i vatten när en grupp människor leker i stadens fontän.
En man med ryggsäck äter en glasstrut.
En kvinna med en kopp och en gäspande man sitter framför Cigar Company-butiken.
En man i blå rock går nerför en trottoar.
En man sitter och läser en tidning i ett rum med en klassisk blå bil.
Leverantörer hökar sina varor på en utomhusmarknad.
Sex flickor i sovrumsgolvet som knäböjer på varandras rygg för att bilda en pyramid.
En man i kostym som pratar med en sittande kvinna.
En medelålders man suger upp solen i en allmän park.
En kvinna som bär vita solglasögon håller i en plastmugg.
En man kastas i luften av en stor grupp som håller i kanterna på en flagga.
En man som hoppar från en byggnad till en fallskärm.
En grupp människor på en gata täckta av skräp och rök.
En gammal man med en cigarett i munnen.
En liten pojke på en kaklad köksgolv håller en röd snabbare.
En kvinna som gör yoga.
Ett äldre par går hand i hand en vacker dag tillsammans nära en livlig gata.
En kvinna visar en liten flicka sin ansiktsmålning med en spegel.
En man som håller sig på toppen av en hoppande häst medan andra står och tittar på honom i en folksamling.
Sportfans firar efter lagets seger.
En man som håller Texas flagga är nästan blåst av fötterna på en gata.
En skadad man ligger på trottoaren med en man som håller i huvudet.
En kvinna i vit topp och jeans promoting för CYFD vid gatan.
En man som fiskar vid en flod.
En liten flicka i rosa kläder tittar rakt fram och håller ett par kikare på en stenig spår.
En man tittar på vad man får i affärerna.
En kvinna med långt hår och en svart skjorta diskar.
En man i vit jacka och hatar fläsk till smörgåsar.
En hindu som sover på golvet.
En man och kvinna som äter äpplen i parken.
En man som bär en stor sombrero går nerför stranden med en kvinna.
Folk samlas för att höra ett tal om den armeniska folkmordet.
En kvinna i mellanöstern pratar in i en mikrofon vid ett protestevenemang.
En man och en kvinna som står med en grupp åskådare.
En flicka i lila tröja ser en pojke dricka ur en flaska.
En kvinna i klänning går under en molnig blå himmel.
En man med hatt sitter på marken med en liten väska.
Den här mannen går nerför gatan med en hand i byxfickan.
En kvinna med rött hår bär en blå klänning och har en stor ryggtatuering.
En man går sin cykel i Kina.
En kvinna i bikini njuter av en dag på stranden vid havet.
Infödda amerikaner i dekorativ klänning verkar fira för en sak.
En liten pojke som sitter framför en affär i ett något utslitet område.
En vagn på väg nerför gatan
En kvinna som ligger framför dörrarna till en grinig, gul, röd och grönfärgad byggnad.
Brunett flicka med ryggsäck redo en färgglad drake.
Barnet sitter på gunga utan en tanke i sitt sinne.
Mannen med många medaljer tittar på tjejen i den gula bikinin.
Flera personer, av vilka en bär en kanindräkt, leker i en offentlig fontän med ballonger i närheten.
Många män i blå uniformer går i formation.
Sex personer sitter på en stenbänk utanför en restaurang och tittar åt olika håll.
Två turister helt enkelt klädda stående framför två bankomater.
En grupp människor i ett "ölträdgårdar", samlades under ett grönt presenningstält.
Flera blå paraplybord där människor äter.
En pojke i röd skjorta som sitter ovanpå en järnvägskorsningsbar.
Indian flicka med sin mamma be eller utföra en ritual
En kvinna går framför en tegelvägg en solig dag.
Turister går på kullerstensgator förbi restaurang.
Två personer cyklar nerför vägen framför en hög, gul och vit byggnad.
Tre män i långa kläder sitter och tillbringar dagen tillsammans.
En kvinna springer fram till en jonglerande man på en lina.
En man i kostym läser tidningen medan han går nerför gatan.
En person går vid en vägg som omger en kyrka.
Två kvinnor sitter på trappan och diskuterar.
En kvinna och några barn står på trottoaren och tittar på en fontän som är frusen.
Ett barn som bär en blå hjälm visas sin cykel från sin far.
Vissa människor tittar på produkter som staplas till försäljning på en marknad.
En röd dubbeldäckare i Europa.
En kvinna i svart jacka och bruna stövlar går på gatan framför en grupp människor.
En flicka i vit skjorta gör en yoga flytta ovanpå en staty.
Hon sänker tänderna till ett välsmakande bett.
Tre personer går nerför en stadsgata.
En man med ett bambubandanna ser ut i fjärran när han håller i en bambufiskespö.
En man med en käpp tittar genom kikaren för att se bergen.
En kvinna i svart t-shirt dammsuger korridoren.
En svart hög hoppare utför ett hopp över en stolpe.
En man med en egyptisk huvudbonad och ingen skjorta på håller upp en docka och ler.
En man med en väska går nerför gatan.
Tre personer bär vitt, medan de går på styltor nerför en väg utomhus.
De är hörlurar i manliga subjekt öron och han har också en iPod.
Flera uniformerade människor står vid uppmärksamheten och en kröns av en officer.
Individer i militärkläder samlas under ett trapphus.
Kvinnan i orange slöja med handen över ansiktet sittandes i en blå stol.
En pojke cyklar med utsikt över en stor vattenförekomst.
En man i solglasögon, en mössa, mörka jeans och en jeansjacka går förbi en båge.
Två kvinnor packar upp något från en låda.
Ett barn som håller i en gul filt tittar i en låda med haklappar och leksaker.
En polis i London som skriver en biljett till en man.
En dam i lila och en dam i blått står med en skåpbil bakom sig.
Fyra unga kvinnor går nerför gatan med stora väskor.
En äldre man i beigejacka står utanför en gammal byggnad och läser en tidning.
Två smala, vackra kvinnor i skumma kläder som går tillsammans.
En man som går nerför en smutsig gata framför en byggnad som har graffiti och affischer på sig.
Med händerna vikta, sitter på en bänk stirrandes på en tom skärm.
En räddningsarbetare tittar ut genom fönstret på ett fordon som rör sig.
En blond sångare framför ett kalejdoskop.
En knasig kvinna sjunger på scenen.
Två man på hingstar utför lassoing en liten svart kalv.
En makeup artist som bär rosa och vitt ansikte färg och garn peruk applicerar ansiktsfärg på ett litet barn.
En ung flicka som står vid kanten av gatan i en vit klänning.
En man i vita shorts är i en park och kastar en frisbee.
Två kvinnor delar paraply.
En ung man, klädd i en svart skjorta med ordet "kärlek" över, jonglera tre gröna bollar.
En kvinna går sin hund på en marknadsplats.
Många människor går längs gatorna framför en stor, grön staty.
Kvinna sjunger på scenen framför backup dansare
Två kvinnor går över en gata, en bär en röd skjorta och rosa hatt, medan den andra bär en randig, vit skjorta och solglasögon
Två damer går tillsammans och har kul.
En kvinna drar upp en motorcykel på ett hjul och utför ett trick.
Den här kvinnan cyklar i underkläderna.
Är äldre person med en blå jacka sittandes på en bänk och äter en glasstrut.
Två tonåringar går nerför gatan med en arm runt en annan.
En skäggig man i svart t-shirt sitter framför ett skrivbord med en dator.
En man slappnar av i skuggan och tittar på stranden.
En äldre skäggig man i någon slags tjusig svart och vit klädsel omgiven av en grupp åskådare.
En kvinna faller genom luften.
Fem pojkar som två har en skateboard framför statyn.
Kvinnan på en marknad får lite frukt.
En kvinna med mikrofon står bredvid en man som använder en Apple-dator.
En man som ser en dam korsa gatan.
En äldre afroamerikansk man som har lotter på en gata.
En man står i en folkmassa och håller upp ett tecken.
En massa människor är med sina cyklar som bara bär sina underkläder.
En dam med ljust orange hår som går i en folkmassa.
Två gamla människor sitter i stolar på trottoaren framför husen.
En ung rödhårig flicka avslutar sin lunch.
Två äldre kvinnor undersöker en utställningslåda med föremål till salu.
Foto taget inifrån en restaurang av människor på gatan.
Dessa unga damer sitter bekvämt diskuterar sin mat eller talar om kvinnan.
En man med en gul skjorta på stirrar i fjärran
En äldre herre som håller en burk kokain och en ung pojke är på något slags marknadsevenemang och tittar på något till salu.
En ung dam som sitter utanför ett sportevenemang och tittar på sin telefon.
En man och två kvinnor provar olika födoämnen.
Flera äldre personer står framför ett matbås.
En kvinna på en kiosk dekorera kopp kakor medan åskådare uppmärksamt observera tekniken.
Kvinnor lagar stekt mat på en utomhusmarknad.
Två personer tittar på en uppvisning av flaskor.
En man med blå handskar lagar mat under ett tält.
Två kvinnor står tillsammans bland en skara människor som äter lite mat.
En man i gul skjorta som går och dricker en öl.
Kvinnan i lila tröja talar medan hennes vän i grön tröja lyssnar.
En svart man med rosa skjorta sitter på en busshållplats och röker en cigarett.
En grupp unga damer med skyltar är på gatan och protesterar mot oljeutsläpp.
Folk på en gata delar sina åsikter om olja.
Hemlösa människor sover på gatan framför en affär.
En massa människor på en karneval.
En cyklist i orange shorts och grön ryggsäck som passerar genom en livlig gata.
Två små barn leker i smutsen med spadar.
En ovanligt klädd man med sin enhjuling och sin ovanligt klädda partner.
En asiatisk kvinna äter mat med andra människor.
Två killar klättrar upp i ett träd för en bättre utsikt över vattnet.
En person hoppar i luften, med snö på marken och massor av träd i bakgrunden.
Två kvinnor pratar i ett bås som är fullt av hattar.
Två kvinnor besöker ett vin provbord.
Folk står i kö för öl och curry.
Det högra hörnet är böjt på höger sida, det blå vitt och grönt.
En ung man säljer isglass och läsk med en tröja på höfterna.
En grupp människor samlas på gatan.
En grupp människor står runt ett matbord medan två personer serverar sig själva.
En äldre man arbetar för att sälja bröd till en äldre kvinna.
En ung man med vit hatt och svart skjorta blandar fruktdrycker för människor.
Människor står och går runt framför ett shoppingområde.
En kvinna sträcker sig efter något i sin väska när de står framför ett matstånd.
Band som spelar utomhus inför en grupp människor.
En utländsk man i svart och brun hatt står stilla mitt på trottoaren.
En kvinna i vit skjorta som går på trottoaren.
En grupp män som bär hattar och skyddsvästar står på en stor metallstruktur.
Bronislaw Komorowskis kampanjskylt svävar över en McDonald's.
En grupp människor i vita sportkläder samlas tillsammans medan en av dem utför en dans.
Åskådare tittar på en ung pojke klädd i traditionella kläder medan de går längs en väg.
En kvinna i lila klänning, som håller en öl, går i en stor skara människor.
En brandman med en brinnande byggnad i bakgrunden.
En man i blå mössa som gör sig redo att fotografera en scen.
En grupp brandmän går nerför en gata.
Människorna är på stranden och tittar på havets skönhet med hjälp av ett teleskop.
En brandman som går under det röda repet.
En grupp brandmän rör sig i ett begränsat område.
Några brandmän har blockerat gatan och folk tittar bakom bandet.
En kvinna som bär en lila klänning med en blå ryggsäck fixar håret samtidigt som hon bär solglasögon
En man går vid en vägg täckt av graffiti.
Gamlingen med svarta Barret och glasögon tittar på en tidning när han går förbi en gammal byggnad.
Flera nyhetsmedarbetare håller ut mikrofoner till två män.
En man som bär brandmansrock och hatt tittar nerför en öppning.
En brandman är utanför stan.
En man som går i staden bredvid en grupp duvor.
En brandman är på gatan och tittar ner.
En grupp människor rider skotrar och motorcyklar på en gata.
2 personer tillagar kaffe på en butik.
Ett antal personer som står på trottoaren längs med ytterdörrarna till en transitbuss
Asiater som bär hjälm och väntar på att få köpa mat.
Brandmännen försöker få isär bilen för att nåt hemskt har hänt.
En kvinna står utanför en byggnad och pratar på sin mobil.
4 personer kanot nerför en flod i en gammal kanot som ligger lågt i vattnet.
Två kvinnor, en man, och två hundar upptar ett gathörn.
En man som går nerför piren och kliar sig i ryggen med en båt som seglar i bakgrunden när solen går ner över vattnet.
En mörkhårig man i en brun t-shirt som går på gatan.
En man i kostym lutar sig tillbaka på en bänk i en busshållplats.
Sju barn runt en vagn som är full av tegel
En man som bär sandal, går nerför en skogsväg mot vatten och bär en handduk och en strandväska.
En man kollar en vägg.
Två män och en kvinnlig vandrare, alla klädda i t-shirts och shorts, poserar framför en spårkarta i snön.
En kvinna som läser i parken med skorna av.
Folk tittade på konst som representerar en osynlig man gjord av en svart kostym och hade ett regnbågsfärgat paraply.
Två personer sitter och njuter av en del drycker.
En ung pojke i en blå jacka som står på ett hörn framför THEFACESHOP.
En man i kostym står i en grupp människor.
En dam står och tittar på alla kläder på marken.
En man har sin handdator och tittar på en lista över flygningar på flygplatsen.
En man står i sanden och kastar en bönsäck i ett hål.
Två män bär västar håller rökiga facklor
Min, låt oss titta på när den vita och röda bilen toppar över.
Arbetare tar fram en mall från en lastbil.
En kvinna i röd skjorta och denimkjol fotograferar en skulptur som omges av byggnadsstaket.
En man som städar ett föremål i fontänen.
En man i grön skjorta och blå jeans står på en korsning mittemot en stor byggnad.
En kvinna och ett barn är på väg att spela tennis.
Två män i röda skjortor som bär en glasruta över en gatukorsning.
Folk går genom ett köpcentrum.
En man som bär förkläde lagar mat i ett kök.
En man med orange overall ger en presentation på ett utomhusevenemang.
Ett litet barn klädd i gula danser bland en grupp människor samlades utanför.
Hunden återvänder med jägarens fågel.
En äldre kvinna som bär en grön klänning håller en käpp och går längs en planterad gångväg.
En Lakers fan fest med människor som håller gula Lakers flaggor.
En kvinna håller en man vid kragen på trottoarkanten när en buss närmar sig på gatan.
En mor bär sitt barn genom en marknad på ryggen.
En ung man som bär en vit skjorta med en karaktär som beskrivs mycket mörkt.
En muslimsk kvinna ligger i öknens öde sand.
En man och en kvinna går framför en vit pickup och en grå bil.
Gamlingen underhåller sin familj genom att spela dragspel
En man sitter utanför med sin resväska öppen och spelar dragspel.
En man i jeans som drar i en resväska.
En skara människor sitter i stolar utomhus, med en stadsscen och en bro i den omedelbara bakgrunden.
Folk äter under ett randigt rött och vitt överhäng.
Två personer handlar i en stormarknad med internationella flaggor ovanför huvudet.
En vy över folk som tittar på en butiksgång.
En gammal kvinna i blå tröja och svart klänning sitter på en bänk.
En kvinna i svart och högklackat med röd väska går.
En kvinna med blå jacka äter lunch med en vän.
En gammal dam som håller i en kamera.
En brunhyad man i en grön tröja med huva och blå jeans bär hörlurar anslutna till en handhållen enhet.
Två små flickor med rosa kläder dansar tillsammans.
Utrustade ryttare rider sadlade och betslade hästar går genom höga gröna gräs.
Människor tycker om att handla färska produkter på en bondemarknad.
En kvinna köper kött på en stormarknad.
Många kunder surfar efter produkter på en marknad.
Två personer som jobbar i en bagelbutik, som firar 20-års jubileum.
Vissa människor tittar på val i en inomhus matplan.
Arbetare i ett kök på en restaurang syns genom ett skyltfönster.
En man som lagar mat i ett kök.
En kvinna tittar på färskt kött och skaldjur i en deli i en livsmedelsbutik.
Fyra personer surfar på en marknad.
Köpmän som går nerför en ö i en livsmedelsbutik.
Folk handlar varor i ett fruktstånd.
Många människor genomsöker den öppna marknaden för internationella livsmedelslager.
Två kvinnor och ett barn i en affär.
En långhårig man i shorts som går nerför gatan med en käpp.
En man som griper tag i ett vitt pappersark sitter bredvid hamnen.
En man i röd skjorta och shorts går längs trottoaren förbi ett Pizza Inn.
Många människor dansar på en stor sammankomst på natten.
En liten flicka med blont hår klädd i en svart tank topp och en kjol vattna utomhus växter med en slang.
En ung pojke hoppar från en dykbräda.
En liten grupp människor under ett träd med en vit pick-up lastbil i bakgrunden.
En gata fylld med människor som går och cyklar.
En grupp barn som poserar med sina intyg.
En mängd olika passagerare åker en turbuss nerför gatan.
Flera personer går längs en gata i tennisskor och shorts.
Många människor med paraplyer går i regnet.
Vackert klädd kvinna posera för bilder eller stå och prata, medan förbipasserande promenader vid en fontän.
Ett par omfamnar på en livlig gata.
En kvinna ringer en mobiltelefon medan hon går förbi en butik med en reflektion i fönstret.
Kvinnlig joggare löper längs en flod i en stad.
En man som bär hjälm kör en ljusröd motorcykel i trafiken.
En kvinna läser en bok och en man passerar tiden på tunnelbanan.
En orientalisk kvinna som tvättar något i ett badkar med vatten och tvål.
Två vänner njuter av glass på en trevlig dag.
En gråhårig man med glasögon och klädd i randiga skjortaffärer för frukt
En person placerar bilmattor på marken.
En ljusbrun valp som bär en munkorg står upprätt mot en kvinna med röda naglar.
En full papperskorg med graffiti på.
En man spelar trummor på en stadsgata.
Jordbrukarna ställer upp sig och tar hand om sin boskap.
En person i svarta shorts, medan skjorta och vit hatt, ler i en publik när hon håller sin cykel.
Folk går genom en fullsatt marknad.
En person håller ett gäng ballonger, varav många är av SvampBob Squarepants.
En man med röd skjorta som städar grillen.
En svart kille med dreadlocks dansar tillsammans med andra människor.
En man som serverar öl från kranen när kvinnan väntar.
Ett rockband som uppträder på en scen en gitarrist, sångare och en trummis
En man som spelar ett instrument på scenen.
En mörkhårig man med randig skjorta som sitter ute med en fruktvagn för att göra drycker.
Ett barn i grön skjorta befinner sig i ett trångt klassrum.
En man i jacka och hatt tar en paus från sin bekantskap och sin drink för en tummar upp
Tjej i hatt och solglasögon tittar på något i fjärran.
En svart hund framför ett träd som hoppar mot en röd frisbee.
En tjej jobbar med sin tränare på en gymnastikbar.
En flicka i en rosa solklänning skjuter en skoter förbi en rad orange byggfat.
Två unga vuxna som korsar gatan med hjälp av en trottoar.
En äldre man sitter på en bänk framför ett gräsbevuxen område.
En person går upp för yttertrappan mellan två byggnader.
En räddningsarbetare som gör sig redo att bända upp en bil som har vänt över
En man i ett fordon pekar på något.
En liten flicka, klädd i rosa och vitt med blommor i håret, står utanför och rör vid hennes bröst.
En man sitter och läser en bok.
Tre män sitter ovanpå en grön tank.
En man på gatan stirrar på en vagn.
Två män sitter på lägerstolar medan de läser eller studerar.
En person som samlar blommor i en silverskål.
Flygfoto över fotgängare som går på trottoaren på en gata i en livlig del av staden med träd i median.
En person som jobbar på en matvagn.
Det är en man som fiskar på en bro.
Färgglada tecken med asiatiska karaktärer lyser upp en gränd på natten.
En grupp människor protesterar med tecken som säger: "Sluta döda i Iran."
De dansar på gatorna topless.
Mannen i den gröna rutiga skjortan äter något.
En livlig grupp civila är i staden.
Ett band spelar på en scen med lila spotlights.
En man arbetar med ett byggprojekt utanför en byggnad.
En man med blå hatt står bredvid några cyklar och en massa människor.
Folk tittar på en fotbollsmatch vid det lokala vattenhålet.
Folk sitter utanför ett café och äter och dricker.
En kvinna är i en spritbutik.
Folk sitter på piren vid kanten av vattnet.
Matförsäljaren går sin vagn med mat längs en väg.
Folk sitter på bänkar på en trottoar omgiven av träd med utsikt över stadens byggnader.
En dörr större står vid en öppen dörr till en byggnad.
Folk går längs en tegelstensgator som är fodrad med affärer under en molnig himmel.
En grupp bargäster njuter av fotbollsmatchen.
Cyklister rider genom en skog medan åskådare hejar.
De cyklar på gatorna.
En biker i vita kläder tar händerna från styret mitt på en skogsväg.
En grupp cyklister cyklar nerför en väg.
Åtta personer är på en rulltrappa som går upp eller ner.
Folk går längs trottoaren en kall dag.
Två kvinnor i bikini toppar och shorts går vid en sjö med två män.
En man i röd skjorta tittar på ett fallet träd.
4 medlemmar i ett band spelar tillsammans utanför på en trottoar.
Gatumusiker i röda dräkter som spelar på trottoaren.
En kvinna går sin väg på en trägång genom ett fält av gyllene växter.
En äldre kvinna går i regnet och håller ett rött paraply över sig.
Asiatisk man med en vit skjorta och grå byxor stående med en mikrofon nära en högtalare.
En man för ett samtal medan en rad individer rör sig bakom honom.
En kvinna håller i kaffe och sin mobiltelefon och verkar leta efter någon.
Ett band spelar musik på scenen.
Ensam person i en kanot, håller i ett rep, njuter av landskapet i de blå bergen och glasigt vatten.
En hona med solglasögon pratar på sin mobil.
En blå båt rör sig nerför en kanal kantad av röda, orange och vita hem.
En kvinna i svart minikjol som cyklar orange.
En folkmassa står på en väg mellan höga byggnader.
En cyklist ringer någon eller kollar hans sms.
En ung man hälsar på sina anhängare innan en stor karatestrid hålls i hans stad
Ett barn med blont lockigt hår som gråter.
Fyra medlemmar i ett band uppträder på scenen.
En man i slips på en gata.
En svart flicka och vit flicka som går hand och hand i ett livligt område i en stad med ett offentligt tåg i bakgrunden.
En jean keps med Tommy Hilfiger-logotypen.
En tonårig blond tjej pratar på mobilen när vinden blåser in håret i hennes ansikte.
En kvinna som bär ryggsäck och glasögon står på en gata.
En kvinna i höga klackar och en kort kjol står mot en tegelvägg på en trottoar.
En man på en bro håller ett blått föremål över rälsen.
En grupp män organiserar en aktivitet på ett gräsfält.
En man övar karate flyttar i silhuett med en bakgrund av en färgstark strand solnedgång.
En man med orange hatt som håller i en pinne pratar med en man som bär solglasögon och har randig skjorta.
En polis lutar sig mot sin motorcykel medan folk tittar.
En grupp människor sitter och stirrar på datorterminaler i ett stort, smalt rum.
Två kvinnor väntar på en tågstation i centrum.
En man i en lång vit skjorta står på gatan.
Ung flicka njuter av sig själv som hon sprejas med en sprinkler
En man som håller i en gitarr med knytnäve i luften.
En tatuerad kvinna bär sina tillhörigheter i en grön ryggsäck.
En man och en kvinna sitter vid ett bord utanför, bredvid en liten blomsterträdgård.
En välklädd man som sträcker ut mat från en kruka i en restaurangmiljö.
En äldre kvinna som knäböjer med en hink inne i ett blått hus.
En äldre man med glasögon håller dörren öppen på en röd minibuss.
En dam och en man sitter på en bänk och pratar och tittar på folk.
En kvinna höjer handen när en buss passerar förbi.
En skallig man som lutar sig mot en byggnad med en ung flicka som hukar sig och håller i en flaska vätska.
Gula banderoller med svart lejonavtryck hänger över några träd i ett solbelyst område.
Kvinnan i brudklänningen står på tegelgången.
En ung man leker i fontänen.
En man i intressanta kläder, bestående av en fjäderhatt, mantel och en utsmyckad käpp, sitter på en bänk utanför en byggnad.
En stor dam och en äldre dam väntar på en busshållplats.
En svart man i blå kostym pratar på en mobiltelefon medan han röker.
En kvinna protesterar mot föroreningar.
Spännande par hoppar så högt de kan medan de njuter av utsikten över bergen.
En man i grå kostym håller tal.
En flicka i en eterisk, blå kostym som håller en dekorerad hulahoop tittar uppmärksamt in i kameran.
Tröjlös man som ligger på en handduk i gräset.
En man, i svarta tajta byxor, sätter sig lutande mot väggen i en vit byggnad.
Ett litet barn som tittar på en leksaksjärnväg.
En kvinna i vit klänning hukar sig i en massa människor.
Tre kvinnor handlar kläder och ett tecken som säger "5 euro".
En ung kvinna smeker den vita kaninen som sitter på benet.
En man går förbi ett porträtt av en man på väggen
En man som bär på ett barn går omkring med en kvinna som håller i ett solparasoll.
En gammal dam bredvid en väggmålning minns att död
En liten flicka klädd i en vit smock med rosa ballonger håller en ljuslykta.
Fyra personer är i vatten och pratar med berg i bakgrunden.
En kvinna som bär en vit klänning och cyklar.
En kvinna i vit klänning som går förbi ett östeuropeiskt tecken.
Två knappt klädda kvinnor kysser varandra i en skara människor.
Två asiatiska män i vita dräkter ber.
Flera män sitter utanför på tegelkanter byggda runt höga träd.
Ett orientaliskt par går förbi en korridor i ett konstmuseum.
En äldre grönsaksförsäljare på utomhusmarknaden sitter med sina varor och läser en tidning.
Tre vikingar går på strandpromenaden.
En ung flicka i svart t-shirt med halsband och armband går nära ett utomhuscafé.
En kvinna poserar med en stor fisk hängande från en krok.
Två män sitter på sina platser med en flicka mellan sig.
Två unga barn spelar något slags spel
En skara människor står utanför ett vitt tåg med flera ingångar.
Våta barn som leker i en parkfontän
Två poliser pratar med två män som har en robot.
En man med en burk går förbi en målning av en byggnadsscen.
En kvinna i bikini ligger på en filt på en brygga över vattnet.
En kvinna i en blacker topp går med sina vänner.
En publik sport färgerna rött, svart och gult på målade ansikten och kläder samtidigt vifta flaggor av samma färg.
En brun och svart hund som skakar om sig själv.
En ung pojke i randig skjorta leker med kvistar på ett gräsfält.
Två lesbiska som mår bra av att bli blöta.
En arbetare i en pizzabutik väntar på att få kunder.
En polis står med armarna korsade.
Omkring 16 män klädda i polisuniformer samlas mitt på en gata.
En manlig magiker som gör ett trick inför en publik.
Tre kvinnor dansar och spelar musik i en grupp.
En grupp människor samlas i en stadsmiljö.
En man med långa dreadlocks stoppas av två män i blå uniformer.
En man ser på medan hans kvinnliga följeslagare täcker hennes ansikte med en servett.
En man i cowboyhatt förbereder korvar på gatan.
Man med glassvagn stående mot en vägg.
En flicka och två pojkar klädda i ljusa etniska kläder går tillsammans.
En grupp om fyra män bär en staty.
En man i gul röd blommig klänning spelar gitarr
En rodeo cowboy rider på en bagatellhäst.
Två män och en kvinna gör yoga i ett vardagsrum.
En kvinna sitter på en bänk framför en elefantutställning på ett museum.
En kvinna i en tank topp och jeans rider sin cykel längs en väg.
En äldre man klipper en yngre man.
Mannen i tanken tvättar ansiktet med vatten från en träskål.
Ett par tittar på en show på en restaurang.
En ung man i korthet, shorts är mitt i en stor publik på sin mobiltelefon.
En man med en vagn full av risrök på gatan.
En kvinna ammar ett barn i vad som verkar vara en marsch.
Människan inspekterar korv inuti en deli.
Ett ungt par är i början av att spela Jenga på ett vardagsrum soffbord.
Polisen med gasmasker knäböjer framför marken.
En man håller sin skjorta i en fontän i en park.
Mörkhårig man sitter på blå stol och tittar på tvättmaskiner.
En liten asiatisk flicka i en blommig klänning står i dörröppningen och håller en nallebjörn och ett mellanmål.
En kvinna håller i ett rött paraply och en fläkt.
En flintskallig man klädd i svart med hjälp av en fläkt gjord av fjädrar, som går nerför gatan.
En man med ett målat ansikte, klädda i damkläder och cyklade.
En man i blå skjorta ställer sig på gatan framför polisen i upploppsdräkt.
Mannen i den vita t-shirten talar på ett podi.
Två män sitter vid en disk och tittar på förstoringsglas samtidigt.
Folk går nerför gatan en solig dag.
En flicka med en lila mohawk och en röd tank övredel pekar och pratar med en skjortlös kille utanför en byggnad.
En man är klädd i en svart prickig hatt och mantel.
Flera figurer i klänningsskjortor och slipsar stirrar ut genom fönstret i en tegelbyggnad.
En man leker med ett barn.
Ett barn är klädd i kostym och håller en treudd.
En blond kvinna korsar gatan i affärskläder.
En man i blå skjorta håller i en skylt och ber om jobb.
Poliser som står utanför en affär.
En kvinna dansar och en man håller i en åra.
En kvinna i lila kjol dansar.
En kvinna som bär en gräskjol och blommor i håret håller en kanna.
En äldre man som plockar blommor.
En man sitter framför en fruktvagn och vinkar åt någon.
En kvinna skuggar sig från solen med sitt paraply.
Två män och en kvinna sitter på en bänk, nära vatten.
En blomsterflicka poserar i en dörröppning.
Ett äldre par sitter med sin hund på ett grönt fält vid stranden.
En orientalisk dam poserar med svart behå och håller i en näsduk.
Två dansande damer med ryggen mot kameran är i en synkroniserad pose.
En grupp barn vandrar på en stig.
Ett ungt par är utanför bland många andra människor och den unga damen håller i en champagne eller vinflaska.
Tre vuxna odlar framför ett metallstängsel.
En man står på en livlig trottoar med en Brasilienskjorta och viftar med en Brasilienflagga.
Tre gamla män sitter ner och pratar.
Solskenet som lyser in utifrån ger en vanlig indisk kvinna ett ögonblicks klarhet.
En kvinna kramar en skjortlös man.
Två mörkhåriga kvinnor sitter på gråa steg bakom ett grått staket.
Ett par går sin Dachshund förbi en vägg med graffiti på.
En ung flicka i blå skjorta och denimshorts, som drar i ett rep och står i en grop av lera.
En ung flicka som leker på en lekplats.
Medan han är i Schweiz väntar en man i en blå tröja för länge och tar en öl.
Människor som står nära ett stort metalliserat föremål som speglar en stads skyline.
En man och en kvinna knäböjer utanför, ritar ett stort porträtt på betongen av en kvinna som håller ett barn
En person i en blå skjorta sover i ett gammalt monument.
Två kvinnor deltar i en drakdans.
Många människor samlades utanför, satt på bänkar och i gräs.
Två unga män som bär solglasögon och vita poloskjortor står utomhus och tittar på tidningar.
En skjortlös man läser sportavsnittet i en tidning.
En man går en hund på en tom väg.
En gata full av affärer.
Två poliser förhör en sittande man framför ett tunnelbanetåg.
En man som sticker en metallstav i en flod av lava.
Tjejen som står längst bak i husvagnen och ler när hon rör på höet.
Akutmedicinare arbetar för att hjälpa en man.
En kvinna som går två hundar framför en vägg med en strand dragen på den
Ett par stora glasögon som sitter utanför en byggnad.
Ett gathörn med två förbipasserande cyklister och flera fotgängare.
En man bär en väska i sin vänstra hand.
En dam i svart och röd utstyrsel som hoppar över en dam i svart klänning och spelar ett instrument.
En stor folkmassa går stadens gator på natten.
En tjej säljer iste med färska citroner och mynta.
En liten flicka, allt i rosa, ler mot kameran från hennes plats på den vita mattan.
Två ungdomar i shorts och t-shirts spelar basket i en urban utomhusbana.
En man på en stege tvättar en byggnad.
Tjej i tank topp och byxor svänger på en stock sving.
Fotografer tar bilder av saker runt omkring sig.
En man skjuter eld ur munnen medan han håller i en fackla.
En röd skylt som läser "ARRIVO" hänger ovanför en gata.
En liten svart och brun hund hoppar på en stor orange hund.
Kvinna med rött paraply går i en stad.
Blondhårig kvinna i lila tröja äter en chokladglasskon.
Folk som bär baddräkter på en våt yta.
En man med hatt på läser bakom en kvinna i en tung rock.
En ung flicka läser en bok för en annan.
En hemlös man går nerför gatan med en cigarett i munnen.
En man i jeans och en svart skjorta väntar på en parkbänk.
En övergiven väg med en man i röd skjorta som joggar i fjärran.
En ung flicka som bär solglasögon sitter bland en publik.
En afrikansk amerikansk kvinna i en silverfärgad kjol som går.
Det här är en kvinna i gul skjorta som bär en brun handväska.
En ung kvinna spelar ett stränginstrument på en offentlig plats.
En tjej i svart t-shirt och blå jeans som går på vägen.
Tre kvinnor och en man går med ett barn.
En kvinna pratar på sin mobil när hon står nära en tegelvägg.
En kvinna med en orange skjorta som säljer grönsaker på gatan.
Fyra personer bär flytvästar på en motorbåt på stilla vatten.
En tjej i jeansshorts och en blommig blå och grön skjorta lyssnar på sin iPod.
Leverantörer säljer olika varor under stora färgglada paraplyer.
En grupp kraftarbetare på platsen för en bilolycka.
En kvinna i gul skjorta och blå jeansbyxor som går.
Två kvinnor i snygga kläder går nerför gatan.
En kvinna som bär en stor hög med trälådor.
Tre kvinnor ute på gräsmattan i en park område håller motion poserar.
En man med blå jeans ligger ner med huvudet på sin bokväska.
En asiatisk tonåring som bär en vit skjorta med svarta ränder sitter på trappan med ansiktet liggande på handen.
En händelse äger rum utanför.
En grupp människor i en kontorsmiljö som sitter i en cirkel.
En flicka och en pojke som går på stenar.
En man med hatt men ingen skjorta fäster något på en byggnad tak.
Flera videokameror radade upp sig bakom en betongvägg.
En ung kvinna med fåniga gröna glasögon på och en förvirrad blick på ansiktet sitter vid ett bord under ett träd.
Trollkarlen gör ett magiskt trick.
En man hjälper sin dotter med sina skor, vid en simbassäng.
En kvinnlig tennisspelare klädd i vitt med fokus på spelet.
En man med brunt hår som går sin cykel tvärs över gatan.
En flicka står i ett svagt upplyst område.
En kvinna i svart skjorta och blå jeans står på trottoaren
En kvinna med vita solglasögon skrattar.
En dam står bredvid en solfylld byggnad med pelare.
Folk står runt ett bord utanför.
En man som skakar majs medan hans son tittar på TV.
En man med kanadensisk flagga på en fest.
Hon hoppar in i bubbelpoolen med sin ljusrosa badtröja på.
Brandmän reagerar på en motorcykelolycka.
En skallig medelålders man i en tanktopp köper något från en äldre kvinnas bord på en gårdsförsäljning.
En kameraman är på trottoaren och filmar någon klädd i kostym.
Denna Nanny är uppmärksam på de två barn som syns på bilden, och har två andra barnvagnar nära också.
En kvinna som bär motorhuv tittar på en vinflaska.
En ung svart man i grå skjorta som håller upp en skylt på en fullsatt stadsgata.
Vissa människor sitter i en utanför kinesisk restaurang och äter.
En mycket färgstark, full butik i ett köpcentrum, som kallas bris men har festförråd.
Tre nivåer av ett köpcentrum med färgade strängar hängande.
Två kvinnor, en klädd i röd, vit och blå bikini poserar för en bild på en stads gata.
Kvinnor pratar med en äldre kvinna i mycket små kläder.
En stor mängd människor sitter utanför någon form av vattenrelaterade händelse med kanadensiska flaggor.
Människor i röda kanadensiska tröjor sitter på en fontän.
En äldre kvinna i en grå tvådelad outfit jonglerar tennisbollar.
Människor som alla är ute i kanadensiska färger äter mat på en kanadensisk festival.
Ett ungt barn i orange t-shirt rider i en barnvagn.
En rödhårig flicka äter ett potatischips.
Det går människor längs en trottoar i en japansk stad.
En grupp tar sig an ett område som är dekorerat i asiatisk kultur.
Flera personer går på en trottoar bredvid en hög struktur med en väggmålad på den.
Observatörer stirrar på ett stort julgran på trottoaren.
Folk går nära en trottoarvisning som ligger framför en butik.
Tre barn står utanför med en fågel som flyger förbi.
En kvinna i en prickig skjorta väntar på ett säkert ögonblick att korsa gatan.
Män och kvinnor står i ett gathörn.
Foto av en gata i Kinatown delen av USA stad
Några män och barn går på en orientalisk sidogata.
Folk väntar på en korsning bredvid ett trafikljus.
Två personer går i ett storstadsområde nära höga byggnader med skyltar.
Ekonomin hackar och påverkar Kina.
Folk går in i en affär.
En man med shorts tittar på sin mobil medan en kvinna går utanför en liten byggnad.
Tunnelbanetunneln med folk runt omkring
En orientalisk man som bär en budbärarväska och cyklar på en orientalisk gata.
En man som siktar en kamera på något ovanför en gata.
En man som håller kameran över huvudet tar en bild, medan andra sitter i närheten.
Flera asiatiska människor på gatan tittar upp och håller kameror för att spela in något.
En dam som bär jeans och en tanktopp och bär ett paraply rider sin cykel över en gata.
Folk går på en trottoar bredvid en trappa
En asiatisk man med blå skjorta och bruna byxor kör motorcykel.
En äldre man går i en park med två glasstrutar.
En filmaffisch av en man i blått som håller en kvinna i rött utanför en teater
Kinesiskt nyår firas i köpcentret.
En ung flicka i färgglada leggings bär en färgglad flagga i en parad.
Folk spelar fotboll på gräset.
Två ungdomar står i dörröppningen till ett rum fyllt med rosa, vita och röda ballonger.
En man och en kvinna i kostym går framför en vägg.
2 rader kvinna går mot varandra på trottoaren utanför en butik med en pojke 50 % skylt på den gyllene inramade fönster.
En man, klädd i svart hatt, snidar en design i trä.
En scen på en gata, där den ena har shoppingväskor och den andra frågar efter vägen.
En man sitter på marken under ett tecken.
Två flickor går nerför gatan och tittar på föremål i skyltfönster.
En ung man i blått bär utrustning över en gata.
En dam sitter i en stol, framför en graffititäckt vägg med en vagn full av väskor.
En gammal man som sitter i en parkerad gatustädare öppnar dörren.
En pojke klädd i blå racing coveralls sitter på en fotbollsboll på en betong picknick bänk.
En man på en lantlig plats som arbetar för att rentvå ett får.
En äldre man står på en stege och sköter löven på ett träd.
Två clowner står bredvid en kvinna.
En ung pojke på en sele klättrar upp för ett stenblock.
Två svarta kvinnor som går i New York.
Kvinnan i den vita klänningen ser väldigt obekväm ut i de hektiska omgivningarna.
En gammal kvinna som sitter på en bänk.
En man bär sin jacka när han går förbi någon utsmyckad graffiti på en vägg.
En cyklist kör förbi en byggnad täckt av graffiti.
Ett klassiskt propellerdrivet flygplan flyger på avstånd när två män leker med ett fjärrstyrt leksaksflygplan i ett fält i förgrunden.
Två äldre män ute på ett fält på väg att flyga ett leksakskrigsplan.
Det finns 6 unga män som spelar basket i blå och vita uniformer, medan folk tittar på från läktarna.
En man som jobbar på ett litet modellflygplan.
En man i en blå vindjacka leker med sitt gula fjärrstyrda flygplan.
Gammal man i jeans och rutig skjorta hjälper en modell flygplan flyga.
Medan de skyddar sina ögon, väntar tålmodiga åskådare på solförmörkelsens ankomst.
Två äldre människor står nära ett modellflygplan i ett fält.
En person i ett stort fält leker med ett modellflygplan.
Tre män i ett fält med modellflygplan.
Killen med solglasögon och hatt sjunger in i en mikrofon.
Ung man på en soffa fingrar en stor elektronisk tangentbord enhet.
En flicka i en grön tanktopp matar duvor.
En man går längs sidan en ung flicka som cyklar.
Flera personer dricker och pratar vid ett utomhusbord på en restaurang.
En man som står med ett glas i handen och en vit hatt.
En äldre man går i ett stort gräsområde med ett litet plan i bakgrunden som är på väg att landa.
Vackra färgstarka kostymer som visas i en indisk parad.
Folk går och det finns en kvinna klädd i svart klänning och svart huva och fåglar är på trappan.
Någon sitter stilla på en orange motorcykel på en crosswalk, bär en svart väst och hjälm.
Tre barn går förbi ett parkeringsgarage, en av dem är på en cykel.
Folk som står på en tågstation och väntar på tåget.
En kvinna som bär en vit klänning och en blommig handväska har en stor fetatuering på ryggen.
En vit hund simmar med en pinne.
En vit man som bär denim coveralls och en vit baseball keps ser två män som sitter på hinkar spela musik framför en butik som säljer peruker.
En man och en kvinna hoppar upp i luften ivrigt på en träbro.
Här är en bild av en man som går ensam vid oceanpiren.
Flera kvinnor klädda i burkas och ett barn i en orange skjorta ute på en offentlig plats.
Två tonåringar på en skatepark mitt i regnet.
Folk går, sitter och står utanför ett varuhus.
En man fokuserade på att spela sin akustiska gitarr på en trottoar.
Två unga kvinnor går nerför gatan en varm dag.
Två honor (i blå respektive ljus orange skjorta) tar en promenad.
En man går från en bro framför en stor orange byggnad.
En liten flicka i en blå topp och mössa som sitter i gräset och slickar på fingrarna.
En kvinna i eklektisk dräkt drar på en annan kvinnas hand.
Många människor tycks ta en bild.
En grupp personer i badkläder står på ett fält täckt av tält.
En grupp ungdomar tar en löjlig bild framför en kamelstaty utanför.
Unge pojke som håller solglasögon och bär baddräkt.
En grupp män som uppträder som ett band utanför en byggnad.
En man som står på en grön båt.
Tre kvinnor går nerför en tunnel medan en sittande man tittar på dem.
En kvinna läser en bok på tunnelbanan.
Två personer står medan andra går eller rusar förbi.
En man och en kvinna sitter på trappan utomhus och pratar.
Tre kinesiska kvinnor och en man dansar för en publik.
Återuppträdande av gammaldags valsning med kostymer - 3 par
En ung pojke med blont hår och blå ögon står mitt i en lastbil säng med vattenmeloner medan familjemedlemmar står i bakgrunden.
Folk går tillsammans på en gata.
Fem personer, tre kvinnor och två män, utför en dans i period kostym bär utanför.
En kvinna som sitter på några trappsteg röker en cigarett när hon kommer åt sin laptop.
Ett litet barn i röda byxor och en svart kimino som toppen går.
Två barn leker på en stenstrand vid vattnet
Två personer åker motorcykel på en väg framför affärerna.
Två kvinnor går över en gata framför en motorcykel med två passagerare.
Två personer samtalar på en parkbänk i bakgrunden av en låda memorabilia till salu.
En man och en kvinna i viktorianska kostymer hälsar på varandra.
En svartklädd man tar en tupplur i en grön park.
Män lägger grunden till en byggnad.
Två kvinnor går förbi en byggnad med en stor amerikansk flagga och en man som står i en orange skjorta.
Tre poliser vaktar en affär.
Människor väntar tålmodigt i folkmassan vid brandbilen som de leds av brandmannen.
En publik tittar på fyrverkerier på natten.
En ung pojke i grå t-shirt siktar på en pistol fäst vid en lastbil.
Barn i t-shirts står på ett vått däck.
En man i orange skjorta med en orange stege bredvid en tegelvägg.
En kvinna med rött hår som bär en svart blomklänning knäböjer bredvid ett bagage och tittar på en mobiltelefon.
En stor grupp människor korsar en stadsgata.
Kvinna nära en shoppingvagn som går förbi en anka.
Ett färgat par cyklar med vita väggdäck längs en stadsgata.
Två damer i stora solhatt går nerför gatan.
Många människor sitter sida vid sida på en låg cementvägg som skiljer en gata från butiksfronter.
En kvinna njuter av en drink på en full gata.
Sex män sitter framför en docka, fyra av dem bär blått.
En kvinna utanför solbadar på en filt i bikini.
Tre vänner står vid floden och pratar om gamla historier.
Två kvinnor sitter bredvid en trappa täckt av graffiti.
En man som står och tittar på en datorskärm i en butik.
2 män i vita rockar tittar på i en kinesisk restaurang.
En anka står på en trottoar med en asiatisk kvinna och hennes två söner som går mot den.
En äldre kvinna som sitter i fönstret till en stenbyggnad
En man och en kvinna som bär en hijab stående på en bro när ett fartyg passerar i fjärran.
Två personer talar bredvid en flagga med en ögonbild.
Den äldre busschauffören öppnar dörren för en passagerare som behöver kliva av.
En kvinna i gul skjorta som går förbi en parkeringsplats.
En man i gult är på väg att ta en puff av sin cigarr som hans fru tittar på.
En man tar en bild av en kvinna på en fullsatt gata.
Folk ställer upp sig och väntar på att säkerhetsvakten ska släppa in dem i en händelse.
En man i solglasögon och en rutig skjorta som spelar gitarr.
Två personer, en man och en kvinna, är på en scen i ett band.
Ett ungt par umgås.
Tre unga män ro en luftfylld flotte nerför en betongformad vattenväg.
Ett litet band spelar på en bistro.
Ett brandmanslag sprutar en brinnande och rökande bil med en slang på en korsning.
Folk som ser andra uppträda på scenen.
Tre personer sitter på en buss och gör något annorlunda.
En kvinna med ryggsäck står bredvid en cykel.
En kvinna i svart skjorta blåser en kyss.
En hemlös kvinna sover framför ett altare.
En person bär en grön skjorta medan han sover på trottoaren medan en annan person med svarta byxor sover på trappan.
En stor kvinna som satt framför Beatles berättelseutställning.
En pojke bär en stor väska på huvudet från en skåpbil.
En cowboy faller av en häst på en rodeo.
En man som har en mohawk är på en marknad med en buggy i handen.
En man och en kvinna klädd i ljus orange klädsel
Sex svarta poliser, en vit poliskvinna och en vit polis står utanför.
En far läste en bildbok för sin unga dotter.
En man och en kvinna hoppar från en pire till en sjö.
En man som håller i ett blått bälte som är runt en kvinna i svart morgonrock.
En bensinstation namn m&amp;h med gas priset på $ 2,52.
En blond tjej i en gunga som bär Crocs.
Svart manlig leverantör håller sig sval under sitt vita paraply väntar på kunder.
En man som spelar tangentbord i en tom tunnelbanestation.
En man med vit skjorta och glasögon sitter på marken.
Många kvinnor håller upp en skylt som läser "impeach".
En grupp människor står nära ett träd och spelar instrument.
En man som sitter på en silverstolpe på trottoaren med utsikt över gatan.
Folk går nerför en smal gata som är fodrad med bilar.
En man håller upp en "fria kramar" skylt ovanför huvudet.
En man i en cykel och en man som närmar sig honom pratar med honom och i omgivningen finns det massor av cyklar
En grupp unga vuxna hänger på trottoaren utanför byggnadens ingång.
En grupp asiatiska människor trängs ner på golvet och vilar.
Tre personer använder en hemgjord vagn för att bära vatten från en brunn
Tre män sitter bredvid varandra och tittar åt sidan.
En genomsnittlig man som ser ut att spela gitarr.
En skara kvinnor och män samlas under paraplyer på gatan.
En brunettkvinna målar stor väggmålning på marken.
En man som dammsuger nära ett litet barn i ett mjukt grönt målat rum.
En äldre kvinna tittar på sig själv genom en spegel.
En man i mörk våtdräkt som surfar i ett blått vattenhavet.
Tre pojkar och en mamma i hamnen.
En kvinna id dekorera en pärla att placeras med de andra.
En kvinna övar på att väva på en traditionell vävstol.
En fläckig hund sätter sin mun upp till ett litet barn ansikte som får uppmärksamheten med ett skrynkligt ansikte.
Tonåringen cyklade runt på gården.
En kvinna med hörlurar som håller i en penna och ett papper medan hennes fötter är upphängda på stängsel.
Ett flygskott på en liten pojke som bär på en fotbollsboll.
Två unga damer, en blondin som pratar på mobilen, en brunett som sms:ar, går på sommargatan.
En leende man som bär en fotbollströja bär en hög med videospel.
En pojke spelar på ett djungelgym med en basketboll framför sig.
En man klädd i svarta danser med en kvinna i röd klänning utanför.
En tjej i en blå Hollisterskjorta som går nerför gatan med två påsar för evigt 21.
En ung pojke klättrar upp för ett rep av någon lekplats leksak.
Ett gäng barn och vuxna som leker med olika färgade bollar på en trottoar.
En man spelar trummor i ett marschband.
En man med svart skjorta och blå shorts står i dörröppningen till en butiksfront.
En kvinna som jobbar på sin datorläsning.
En kvinna med mörkt rött hår och en svart hatt som tittar på konst i ett galleri.
Etnisk kvinna bakifrån med blå blomskjorta och rött tyg i flätat hår.
Tre personer på två separata motorcyklar passerar varandra på vad som verkar vara en ras i Asien.
Flera män klädda i blå uniformer marscherar.
En flock människor som går på en gammal gata.
En man i blå joggingplan framför en väggmålning.
En kvinna står längs en gata, gömd vid sitt parasoll.
En skjortlös man vadar i mjukt blått vatten.
En man som cyklar med ett rött och vitt paraply har en bild tagen av en folkmassa.
En turist fotograferar en cyklist med ett paraply.
Två män försöker plöja lite jord bakom en röd motorcykel.
Man med kamera och väska går upp för trappor
En man som bär en gul hjälm med sitt visir upp rider en röd motorcykel.
En man nära en Hawaii-skylt.
Ett japanskt par i kimonos går nerför gatan en regnig dag.
Två asiatiska kvinnor som stod i kimonos, medan de log.
Sju personer, tre sittande och fyra stående, titta på inramad affischkonst i ett galleri.
Folk tittar på en konstutställning.
En rad människor som sitter vid ett barpallsbord och tittar ut ur en glasvägg.
En man med gitarr spelar på gatan för dricks.
En blond tjej med ett instrument på ryggen bär en grå tank topp, grå shorts och slet nylon med en cykel.
En man sitter på en bänk med fötterna på en skateboard.
En flicka går in i poolen medan andra pratar vid sidan om.
En äldre kvinna sitter på trappan till ett stort monument.
En brunett man kysser en gråtande bebis.
En äldre man som sopar gatan.
En kvinna i vit klänning håller ett blått paraply i regnet.
En äldre svart man kör sin cykel längs en trottoar.
En ung man i röd skjorta torkar en vit bil med två tyger.
En grupp människor står i närheten av en byggnad.
En pojke i svart huvtröja sitter på ett steg där det står "moose RVS".
Ett par människor korsar gatan.
En manlig figur som bär en svart skjorta och jeans smetar en gitarr medan han håller i picken med munnen.
Två kvinnor går och viftar flaggor på en nästan tom stad gata.
Runners deltar i ett maraton på stängda stadsgator.
En av brottarna har satt dit motståndaren.
En kvinna får sin cigarett tänd av en man utanför ramen.
Ta en tupplur i parken med vänner.
Barn samlas i ett stort rum för att titta på en organiserad föreställning.
En man och en kvinna med pannband pratar med barn med upplyfta händer.
En grupp människor är på en båt i vattnet.
Tre män sitter ute på stolar med röda säten.
Tre personer går upp för en rulltrappa och en man med en kundvagn kommer nerför rulltrappan.
En kvinna sätter ett band i en liten flickas hår.
Två män och en pojke som står framför en tegelbyggnad tittar upp.
En kvinna med en grön klänning använder en mikrofon.
En grupp av tre skalliga män i rött sitter på ett räcke, röker och pratar.
En kvinna och en man, utanför, njuter av varandras sällskap.
Tre vindsurfare rider vågorna i en hackande vattenförekomst.
Ett barn ligger på en filt under en kvinna.
Flera människor samlas nära ett område med ett träd, massor av cyklar och en del skräp, inklusive gamla däck.
En man i en jacka som skildrar det kanadensiska lönnslövet tittar på en konsert.
En ung asiatisk pojke vinkar runt på natten.
En man målar en stor väggmålning på marken.
Skäggig man som sitter på en bänk bredvid en båt.
Tre kvinnor som bär ärmlösa skjortor är upptagna med något.
Två kvinnor båda bär vita skjortor och svarta byxor, en röker sitter på en fixtur på trottoaren.
En kvinna bär solglasögon och ler.
En stor grupp asiatiska människor poserar för en bild med en stormtrupp
Folk står utanför en liten butik.
Två kvinnor i långa klänningar och huvudbonader köper av en köpman.
En liten pojke tittar på fyrverkerier ute på natten.
En grupp blondhåriga vita killar som ser vilsen ut när de går nerför gatan.
En svart man som bär en vit, kraged knapp är sydd.
En kvinna i svart klänning spelar en ukulele och sjunger medan en hatt bär man följer henne med ett par maracas och en trumma i bakgrunden.
En grupp människor åker på en vagn genom en park.
En man med två barn som bär flytvästar är i en simbassäng.
En glad liten flicka rider på karusellen.
En kvinna går vid en vägg som har en väg, blommor, skunk och en orm målad på den.
Två unga damer sitter i ett vardagsrum med mauve stolar och äter snacks.
En kvinna sitter på en bänk under en sfinxskulptur.
En man som går medan han håller i rosor.
Tre kvinnor står i vattnet bredvid en strand.
En vandrare i grön skjorta tittar in i en dalgång från en brant klippa.
En svart och vit hund leker med en golfboll i sanden.
En fiskare tar sig lite lugn tid att vänta på en fångst.
En man lutar sig mot en staty framför en byggnad.
En blond tjej i lila skjorta och rutiga shorts som leker med en snöreleksak.
En street sprejfärgskonstnär skapar nya verk samtidigt som han visar sin konst.
En man som gick nerför en öde gata, visade från marken.
En man med en kamera engagerar en annan man i samtal på en gata.
Ett barn i en lila och gul dörrvakt gråter.
Två barn leker i vatten som faller från en mosaiktäckt pip.
Mannen trängde in i en telefonkiosk med en rosa skjorta.
Ett japanskt par går förbi en kvinna med en halsduk på huvudet medan hon går nerför gatan.
Ett nyfött barn får hjälp av läkare.
En flicka äter ett grönt äpple utanför medan en annan tittar i fjärran.
Kvinnan i vit skjorta tittar på soffor framför en graffiti täckt byggnad.
En ung man tittar runt ett hörn medan han håller sin telefon i sina händer.
Två personer går nerför en bergsstig.
En oidentifierad krökt gata med tre personer som går bort från kameran.
De två människorna kommer ut från grillbutiken.
En brittisk kunglig vakt på patrull utanför en stenbyggnad.
En asiatisk man flyttar vagnar på trottoaren till sin destination.
Lokala muslimer firar öppnandet av en ny restaurang sponsrad av Channel 1 nyheter.
Folk hänger sig på en karnevalresa.
En grupp människor samlas framför en klädaffär.
En man med mask och olika klädesplagg.
Gamla världens stenhus och gator ser vackra ut i bakgrunden, och svag person kan ses gå.
En kvinna och en äldre man deltar på en åktur tillsammans.
Två män täckta av röd färg eller blod på en livlig trottoar.
Folk klädda som zombier paraderar.
Fem personer låtsas vara zombier och ett spädbarn.
Folk går på en gata.
En kvinna i en kort röd klänning och kostym vingar går i en offentlig fontän.
En dam bär en rosa cowboyhatt.
En kvinna med röd hårslips och svart prick som håller en flaska vatten.
En kvinna som bär en flerfärgad solklänning går med en man som bär en svart t-shirt och har nyanser.
En gammal kvinna vaggar sin handrullade cigarett när hon röker.
En ung kvinna som bär randig rockklättring.
Personen med den röda långärmade skjortan klättrar upp för en sten i snön.
Asiatisk kvinna i lila står där på en utländsk plats.
En kvinna i shorts och knähöga strumpor går nerför trottoaren.
En man går med en käpp.
En cykelpolis eller säkerhetsvakt rider framför ett hus.
Folk beter sig som en zombie.
Man med stjärna tatuering bär svart t-shirt och shorts beundra konst visas utanför.
Mannen med den röda slipsen gör ansikten.
En man i lila skjorta och en svart hatt tar en bild med en gul digital kamera
En man tar en bild av en fågel i vattnet.
En man i vit skjorta och mörka byxor går nerför en gata.
Två män samtalar tillsammans klädda i traditionella kläder.
Asiatisk man i blå asiatisk dräkt som dansar inför asiatiska musiker i blått.
En man med skägg i vit rock som ska äta något.
En man och en kvinna i sjal sätter sig framför en vattensamling.
En dam som blir arresterad av en kvinnlig polis.
En man och kvinna som sitter utanför en affär bredvid en tom väg.
Några människor vandrar runt i en gammal, söndersmulad del av en stad.
En man och kvinna i en salong går in i en hall.
En kvinna står framför en byggnad.
En äldre kvinna i en kimono lyssnar på något med hörlurar.
Två barn med svart hår som äter med ätpinnar.
En pojke och flicka leker i en fontän.
En man står på en bro och jobbar.
En vit man ses i en swimmingpool flytande ovanför många flytande modeller.
En kvinna i stövlar står under sitt paraply och pratar i telefon.
En svart man står med ett ben på en kort vägg och pratar på sin mobil.
En tjej i svart skjorta tittar på en kemisk reaktion.
En grupp barn står utanför på en gata.
En kvinna som plockar igenom sitt barns hår.
En man i röd hatt bär en svart övernattningsväska, medan en annan i en cowboyhatt följer honom.
Kvinnan går upp för trappan i ett konstgalleri.
En kvinna står i en publik med en grön skjorta, rosa ryggsäck och en mexikansk flagga fäst vid väskan.
En pojke som håller i en svamp och diskar.
En man står bakom en svart grind.
En kvinna med lila hår är bredvid en man.
Högskoleelever som leker i en pöl vatten, mest klädda i rött.
En kvinna som sover på en bänk i baddräkt.
En actionbild av en trummis i en rutig skjorta som går till stan på ett trumset framför en häck.
Två småbarn och en yngre man njuter av sina flaskor.
En man springer nerför ett sandtäckt berg.
En man lutar sig mot en pelare medan han läser en bok
Tre män färdas genom vatten på en motoriserad uppblåsbar flotte.
Kvinna klädd i vitt med ett barn i knät.
En kvinna med halsduk och handskar och med ansiktet målat går förbi.
En mustachioed man spelar dragspel på gatan.
En kvinna beställer glass från en vit man.
Många mörkhåriga människor samlades för något.
En man och en kvinna står ovanpå en struktur.
En äldre man står ensam på en trottoar på natten.
Två män tittar på en våning som håller på att repareras.
Män står runt ett litet tåg utanför.
En hane i en grön randig tank topp skateboard.
En leende byggnadsarbetare som knäböjer.
En pojke i gult kör en skoter på gatan.
En ung kille som spelar för en publik.
En man står på sidan av en gata i en dörröppning.
Två kvinnor i fotboll uniformer spelar fotboll.
En pojke i vit skjorta gör ett trick på sin skateboard på en skateboardpark.
En liten pojke springer på ett stort gräsfält.
Två hundar springer sida vid sida på fältet.
En gammal man sitter på trottoaren och spelar sin akustiska gitarr.
En man i hjälm hoppar på sin cykel.
En man i medeltida rustning rider ovanpå en häst.
En man i en blå tank topp gör pastell konstverk på trottoaren.
En äldre man som går nerför gatan.
En latinoman lutar sig mot en av kylarna i sitt matstånd.
En ung pojke njuter av det svala vattnet.
En ung man i svart skjorta och jeans och som bär en väska till ett musikinstrument går över en gata.
Två kvinnor sitter på en bänk bredvid en bronsstaty.
En man och en kvinna hälsar på varandra på cyklar framför en byggnad.
Skadad dam som sitter och vilar sitt ben på en vandrare
En upprörd flicka sitter på en stock, huvudet i händerna, framför en cykel instängd i ett träd.
Ett formellt klädd par finner ett informellt ögonblick i fontänen.
En grupp människor på en brygga med en båt på andra sidan av kajen.
En förare stirrar ut genom bilfönstret på en katt på gatan.
En man i svart väst viskar i örat på en leende flicka.
En grupp människor står bakom ett stängsel, många fotograferar.
En medelålders haggard ser rödhårig ut i en vit skjorta och silver halsband, lyssnar på en gul telefon.
Folk står och tittar efter nåt.
Kvinna i lång blå klänning lutar sig över nära vit hink på sidan av en gata.
En liten flicka sover på någons axel.
Män i vita kläder bär ett föremål på sina axlar.
Två män jobbar på bygget.
Blond kvinna i en svart kjol business outfit interagerar med en kundservice kvinna.
Damen går genom rader av barn.
En man går framför ett rosa hotell med en gul väska.
En man i en grön tanktopp som håller i magen.
En tonårstjej som har en t-shirt och baddräkt på botten hoppar ner i en vattenförekomst.
En soldat lär barn hur man hanterar en pistol.
Folk samlas på en gata medan en man i hatt sitter i en stol.
En stor shorts gräver i snön en solig eftermiddag.
En man skyfflar snö medan han bär shorts och en rosa skjorta.
Ett litet barn bär rosa står i en dörröppning.
En äldre man, som håller i ett paket, står framför ett tecken som har en flicka med hörlurar.
En man på en skoter och en röd skjorta tittar tillbaka.
Folk är samlade i någon slags affär vid sidan av gatan.
Kvinnor som sitter vid ett bord med en liten eld.
En man i hatt som svänger och ler mot kameran.
En publik vågor röda och gula flaggor.
Två kvinnor i vita toppar står nära en man och en kvinna med bagage på trottoaren.
En fullsatt gata med fotgängare som leds av polis och barriärer.
En man står på baksidan av en sopbil.
Folk går längs gatan med paraplyer.
Barn på kanske, på deras skola, eller kanske, en fältresa.
Tre personer stirrar på en liten målning.
En man som går tvärs över gatan på vägen som säger "håll dig undan".
Två personer är i havet.
Män på en cykel som transporterar olika storlekar av metallskopor.
En stor kran river en konstruktion medan en person som står i närheten på en upphöjd plattform sprutar vatten från en slang.
Fyra kvinnor står med ryggen mot betraktaren, antingen med bikini toppar eller tank toppar på.
En ung vuxen kastar en softball till hemmabas.
Två unga pojkar i uniform äter ris med händerna medan de sitter på marken.
Två kvinnor, en i traditionella mexikanska kläder, hjälper ett barn tvärs över gatan, som en man ser på.
En tjej i blå klänning står bredvid en trästolpe på trottoaren.
Ett barn och en kvinna på gatan i traditionell dräkt.
En man i t-shirt håller ett spädbarn, som sträcker sig efter sitt ansikte.
En barfota kvinna läser en bok längs vattnet.
Två muslimska män med huvudomslag som går i en stad.
En beundrare på en fotbollsmatch bär en lockig röd peruk.
En kvinna med färgstarka kläder går förbi en jeepcherokee bakom ett stängsel.
Två män tittar över vattnet i en liten båt.
En man i overall och handskar ligger under en lastbil.
Folk går nerför en tegelväg kantad av bilar.
En man i rullstol knuffas mot en munk.
En man läser en tidning.
Folk tittar på stranden och en kvinna i en vintopp tar en bild.
Dam i vit klänning med tatuerat ben tittar på väns kamera.
Två män protesterar med skyltar utanför ett Convention Center som har en skylt som säger "eXXXotica Miami Beach".
Två män i jeans går nära en stor stenvägg.
En man som bär vit skjorta och blå jeans går en hund.
En kvinna i vit klänning cyklar.
En trottoarscen med en tjej i vit skjorta som biter i tummen.
En ung man med ryggsäck och blå solglasögon korsar gatan.
En korthårig man i vit skjorta och khakibyxor går fram förbi en svart bil och håller i en vit anteckningsbok.
En man i vit skjorta och slips går tvärs över gatan.
En kvinna med vågigt kort rött hår och glasögon med en solbränd ärmlös skjorta går nerför en gata.
En grupp människor går genom ett köpcentrum eller en tågstation.
En svart man i affärskostym med händer medan en vit man lyssnar.
En man i röd skjorta kysser en annan man.
En man använder sprayfärg på en väggmålning.
En byggnad har flera balkonger med olika växter som växer på sitt staket.
En flicka står på en grusväg när solen går ner.
Fet man och hund sitter framför en staty.
En grupp pojkar i gröna och blå kläder svingar gröna och blå flaggor i luften till en publik som ser ut som de gör.
En cyklist i en cykelbana.
Brandbilen omger en brinnande byggnad på natten och sprutar vatten från olika håll.
Människan testar teleskopet medan lille pojken tittar på, när de står i en minnespark.
En smutscyklist rider uppför en stenig kulle på en motoriserad smutscykel.
Tre kvinnor går på en gata.
En kvinna håller sitt barn utanför ett rött fönster, bredvid en Color TV-skylt.
En person i sandaler är gömd av stora fotbollsbollar.
En kvinna med svart hår och bär allt svart sitter på en sten och tittar i fjärran.
En blå vägskylt är delvis dold av ett närliggande lövverk.
En kvinna med stickad mössa, mörk jacka och brun vågrätt randig skjorta ler när hon åker skridskor med två kvinnor nära bakom sig.
Barn leker i fontäner i en stad.
Dessa två arbetare arbetar på att bygga upp någon form av metallbyggnad.
En man som beundrar landskapet på en okänd plats.
En kvinna i röd rock lämnar en fotobutik.
En man som står i regnet och bär paraply.
Grupper av människor rider nerför en flod i flottar.
En del paddlar i en luftfylld flotte.
Ett barn simmar i en bäck, medan andra väntar med att hoppa från en sten.
En grupp ungdomar seglar och bär flytvästar.
Ett barn och tre katter vilar på en säng.
En gammal man röker genom att sitta i trappan.
En man med randig skjorta har en kamera över axeln.
Två personer går med en hund och använder paraplyer.
En man i en klargrön skjorta och brättemössa sitter med tre andra män på en betonghöjning.
Folk som bär flytvästar sitter i en båtpaddling.
En grupp människor i flytvästar står på ett stort stenblock i bergen.
En man med en blå tjurmask i en skara människor.
En kvinna sätter sig ner för att spela ett casino videospel.
En man som bär glasögon spelar gitarr bakom ett musikstånd.
En kvinna i vit skjorta och grå kjol om hon står under ett vitt paraply.
En person klädd i gul skjorta och kamouflagebyxor går nerför trottoaren.
Ett barn sitter med huvudet på armen i ett rum.
En man som håller i tänger vid en grillfest.
En långhårig man i vit t-shirt och jeans spelar ett tangentbord stående
En lycklig kvinna plockar genom ljusa gröna och vita blommor.
En man i orange rock och sandaler går förbi en blek orange vägg.
En grupp människor tittar genom ett mikroskop.
En kvinna i rött sippar en drink när hon tittar på människorna under henne.
Två unga asiater i shorts väntar vid en trottoarkant.
En kvinna som bär kjol läser en bok på en stenbänk.
Pojke bogserar varmkorvsvagn med man knuffar kärra bakifrån.
En grupp människor går nerför en stad gata utanför byggnader.
En mörk scen är under uppbyggnad.
En man i röd skjorta och en dam i grön skjorta på en silver moped.
En kvinna som bär sandaler knuffar en vagn med grönsaker.
En kvinna som bär en svart klänning lutar sig mot en byggnad som röker en cigarett.
Fyra asiater sitter på en bänk i en byggnad.
En man går nerför trottoaren framför den färgglada byggnaden.
En tonåring i en blå skjorta åker skateboard förbi en Blockbuster-video.
En äldre man som bär en sombrero rider en mobilitetsskoter medan han handlar skor.
En man i svart skjorta står framför ett nödfordon.
En man spelar saxofon medan folk på gatan lyssnar på musiken.
Man står mot blå vägg med skjorta på huvudet
När den blå himlen är täckt av vita, fluffiga moln, står två personer tillsammans nära en sittgrupp med gröna paraplyer.
Många män sitter och äter tillsammans.
Två dansare ger en föreställning på offentlig funktion.
En kvinna går förbi en grupp på tre män.
En grupp äldre män på scenen som ler och klappar händerna.
En man som går över en gräsplätt mitt på en gata.
En stor trasig kvinna i gul skjorta har en rosa axelväska på axeln.
Två män står framför ett sjabbigt grönsaksstånd.
Tre pojkar är i parken och tittar på när barn leker.
En man i gladiatordräkt står på en livlig gata.
En indisk man i hatt sitter och ler.
En kvinna är en blå topp går mitt i en folkmassa.
En kvinna med mörkt hår sitter på stentrappor och ser fram emot.
En äldre man med vit skjorta sitter på trottoaren.
En kvinna i solbränna tar hand om sina varor på marknaden.
En mörkhårig trummis spelar sitt set med entusiasm.
En kvinna som bär en grön Aeropostaleskjorta och ett grönt armband går nerför gatan med huvudet nedåt.
En man i blå skjorta som korsar gatan med udda föremål i händerna.
Fem barn är på en rutschkana, alla klädda i olika färgade kläder.
En man i en matvagn serverar majs.
En man som står bredvid en bil håller upp händerna.
En kvinna med piercing i ansiktet och rött hår.
En ung man i jeans går nerför en trottoar med en hög med papper på huvudet.
Kvinnan går med röda matkassar nerför kullerstensgatan.
En grupp människor äter en måltid i ett trångt utomhusläge.
En äldre man dricker apelsinjuice på ett café.
En person med mörkt hår med en vit tank topp, röda byxor och vita skor går ner för en trottoar med konstverk visas mot en vägg.
En kvinna i lång kjol som går tvärs över gatan.
En liten flicka i rosa skjorta som sitter i en arenabänk.
En familj slappnar av med kallt vatten utanför husbilen.
En man går förbi en byggnad en solig dag.
Ett par fotograferas framför en stor fontän utomhus.
Flera personer står på en cykel rack för att titta på något över blekmedel.
En kvinna blåser bubblor mitt i en folkmassa.
En duva flyger mot en kvinna som är omgiven av en flock duvor.
En grupp elever tittar över en balkong på en senior resa.
En familjecamping med en husbil och sitter runt ett bord.
En trevlig ung dam på en scen dansar och ser mycket vacker.
Flera människor står runt i ett skogsområde, med en fritidsbil i klar utsikt, två äldre män och två barn kan ses, inklusive en ung, leende flicka.
En pojke som står i vattnet håller i en gul fotboll.
En mamma och hennes två barn läste en bok utanför en byggnad med arbetare klädda i orange.
Tre små barn leker i en fontän.
En kvinna i en pool med en ung flicka kastar en fotboll.
Barn och en kvinna leker i en fontän.
Folk står på en fullsatt gata med resväskor.
En grupp äldre män som samlas i vildmarken
En man som bär en färgglad och randig tröja spelar musik på gatan.
Kvinnan i mörk jacka sitter på en bänk.
En kvinnlig sångare och dansare står på scen på en jazzfestival med en vit klänning med blommönster.
En man roddar en båt genom en flod i en stad.
Tre personer står på en betongvägg bredvid havet.
Tre honor hoppar medan de sträcker sig upp i luften.
Männen står på kanten av en riven byggnad.
En man som ler för kameran stående på en parkeringsplats.
En konstnär säljer sina målningar framför ett stort träd i en park
Två kvinnor med Tye färgade bh, flerfärgade halsband och korta denim shorts.
En trött man sover på sin motorcykel på vägkanten.
En man med ryggsäck står längs en trädkantad gata.
En man som poserar med armarna ut medan vikta kläder och lådor ligger på marken.
Folk korsar en gata bredvid en smart bil.
Folk korsar gatan och en man på trottoaren.
En kvinna i blå skjorta och svarta byxor lagar sin vita strumpa.
En man som bär glasögon talar eller sjunger in i en mikrofon.
En lycklig kvinna och en ung vuxen som får sin bild tagen.
En grupp människor som sitter utanför nära väggar som är målade.
En glapp av ungdomar som sitter ovanpå en cementstruktur.
En man i röd, vit och blå shorts fokuserar på något nedan.
En långhårig kille som spelar trummor.
Två kvinnor som bär sjukvårdsuniformer är på en trottoar och den med gula skor hoppar i luften.
En manlig sångare med solglasögon som sjunger för en mikrofon
Medelålders kvinna med vit blus, sitter vid ett bord utanför en restaurang.
En grupp människor samlas på en gata i staden.
En grupp människor väntar längst ner i trappan att två män i kostym går ner.
En kvinna i brun klänning intervjuar två män.
Stora klara björnar sitter på gatan i New York.
Asiater går nerför gatan på en marknad med sina inköp.
En person cyklar i en stad förbi en butik som heter "Kenji".
En kvinna som ligger på ett fält.
Kunder visar objekt i en liten butik som heter "Jump Shop".
Två pojkar cyklar på gatan.
Ett barn och en förälder eller äldre syskon går på en vandring.
Två asiatiska män i svart sitter utanför och pratar.
En ung person i svarta byxor och en brun fedora använder sin mobila enhet på en trottoar.
En pojke bär en svart t-shirt.
En man i vitt pratar med en man i svart när han står på en plattform.
Flera människor väntar på att något ska anlända.
Kvinnan sitter på läktaren i en cowboyhatt och tittar på nån sorts ranchtävling.
Musiker spelar på scenen på Coney Island, NY.
Ett par sitter i varandra och omfamnar varandra när de blickar ut mot floden.
En författare signerar sin bok för ett fan.
Många vuxna och barn äter en måltid i ett offentligt område.
En flicka går förbi ett parkeringsgarage.
Väggkonst och väggmålningar som presenteras på sidan av East Side Hotel proklamerar att de älskar Berlin.
Folk i och utanför båsen vid ett evenemang.
En tjej i röd jacka som spelar gitarr på en mässa eller cirkus.
Ung man med långt mörkt hår spelar gitarr på scenen.
En grupp människor som bär vita kläder och röda stygn går nerför en gata.
En grupp människor sitter bredvid ett koncessionsstånd.
En dotter hjälper sin mamma i köket i den här familjefoto-open.
En gitarrist med långt hår som spelar gitarr på en konsert
En kvinna i hatt går bort från en liten glassförsäljare bil.
Människan går med höga byggnader med reflektioner bakom sig.
En svart kvinna med afro och glasögon som går nerför en gata i Kinatown, pratar i telefon och bär en flerfärgad halsduk.
Två killar som går på vägen.
Ett band spelar musik på scen under blågröna lampor och med röd bakgrund, en vitskjortad DJ som står mitt i scenen.
En person i röd rock spelar elgitarr.
En man som säljer religiösa parafernalia står framför en moské.
Ett par tittar ut i havet från en bro.
Två män med glasögon och stora mustascher med brittiska flaggor i bakgrunden.
Det här är ett sånt ställe som du kanske ser nästan vad som helst.
Två kvinnor som bär matchande kjolar med Union Jacks tryckta på dem går genom en mässa.
En kille som spelar gitarr på en scen ler.
En kvinna som ligger i ett gräsfält och tar ett foto med sin kamera.
En kvinna som bär en grön t-shirt lutar sig mot en vit kolumn.
En kvinna med rödhårigt överdrag står med en man som bär en skjorta med ränder på.
En svart man i en tanktopp vilar.
Två kvinnor med paraplyer går mellan två bilar när de korsar gatan.
Hunden sover utomhus på den cementerade gatan i asiatiska landet.
En gråhårig dam står bredvid en grönsaksutställning på marknaden.
Tre glada små flickor poserar för ett fotografi.
En man sitter i passagerarsätet på en röd trehjulig rickshaw.
En man i hatt och en orange jacka står bredvid en plast inslagen kvinnlig skyltdocka.
En ung flicka leker bredvid en brandpost som sprutar vatten.
En man och en kvinna klädd i grönt stå förutom en pelare.
En grupp människor som består av 6 personer väntar någonstans medan fyra av dem pratar med varandra.
En hora i ett gathörn.
En kvinna i baddräkt och shorts går nerför gatan i svart hatt och solglasögon.
Man med tillbaka till kameran tittar ut över en skog.
En kvinna i kjol pratar i telefon utanför en restaurang.
Två män sitter tillsammans med en kalender på väggen bakom dem.
En man i rutig skjorta och vita sandaler sover medan han läser tidningen.
En man som tittar bort från kameran sittandes på en vattenfärgad pall.
En familj med små barn med resväskor går nerför ett stenlagt område.
En man och barn drar väskor bakom dem nära en stor glob.
Två uniformerade män pratar medan de står på en väg.
Person som står på trottoaren bredvid högen med sopor.
Två människor sitter runt ett träd och en man poserar vid trädet.
En tjej i jeans sitter på sten och får sin bild tagen.
En man säljer färsk frukt på marknaden.
En stor dam i gul skjorta som håller upp en skylt på spanska.
En gentleman med röd skjorta, glasögon och grått hår står i ett rum fullt av sittande människor.
Tre personer sitter vid ett bord tillsammans.
En kvinna i grön skjorta och svart hjälm kämpar med en man i jeans och en ljusblå skjorta.
En skara människor som väntar längs sidan av en byggnad.
En man i vit skjorta spelar cello bredvid en svart kvinna som spelar harpa.
När du kämpar för att arbeta på byggnadsställningar i fuktigt väder.
Mannen med cykeln väntar på att bilen ska passera så att han kan korsa gatan.
En man i svart svit som pratar podi.
Tre män sitter på en sten avsats, och en har en cigarett i munnen.
En ung man bär flaggor utanför en byggnad
En man som kör en vagn och två hästar går längs gatan
En grupp pojkar som spelar fotboll.
En gammal man, bakom honom på glas, finns många politiska annonser.
En kvinna i blå klänning går på en trottoar.
En kvinna i en blå randig skjorta pratar med någon på gatan.
En kvinna i svart går förbi ett varuhusfönster.
En man i kostym håller en amerikansk flagga bredvid en vit skärm med en logotyp på.
Par som håller händerna på trottoaren framför huset.
En skara människor i vita och röda kläder marscherar genom en röd dörröppning in i en vit gränd, två män med koppar som tittar på till höger.
Två äldre män väntar på att gå över gatan.
En skara människor protesterar med en man i förgrunden.
En man som bär vit skjorta kör en cykel nerför trottoaren.
En ung flicka med en kort röd klänning ringer ett telefonsamtal medan hon håller i en klarblå väska.
Sittande kille som hanterar en häftapparat medan en annan kille tittar på.
Två honor och en hane sitter vid ett bord och äter.
En del asiater samlas för ett evenemang i ett gymnasium.
Två kvinnor, som båda bär svarta skjortor, äter.
Personer med gula skjortor deltar i en konsert.
Många elever som väntar på transport i väntrummet tar bilder på varandra innan de återvänder hem.
Barn som spelar i ett hopphus med ett SvampBob tema.
En grupp barn som sitter vid ett bord håller ett vitt papper.
Två flickor står bakom en annan flicka.
En man med randig skjorta ler och pekar när han har halsband.
Tre personer sitter på bänkar och tittar på folk i parken.
Några cykelcyklister rider på en stig genom en stad.
En skjortlös man med fasor som leker med batonger.
En Boston Celtics fan som äter lunch innan matchen mellan Boston och Lakers.
En skallig man med skägg spelar dragspel framför gröna dörrar
En man och en skrattande kvinna sitter vid ett blått bord med en styrofoamlåda på.
En kvinna som tejpar en papperslapp på en bräda.
Två män sitter på en bänk där en har huvudet i knät och en stor gul väska bredvid honom.
Man med ryggsäck hängande en skylt på en stolpe i en lobby.
En pojke som pekar på nummer ett och ger nummer ett med fingret.
En man och en kvinna som står bredvid varandra skakar hand.
Fyra unga asiatiska kvinnor står utanför vid en tom kartong och använder sugrör för att dricka ur gula koppar.
De tre människorna pratar med varandra.
Unga barn som visar ett spel de spelar i sitt land.
En man och ett barn köper glass av en man med en handskjuten glassbil.
Två män och en kvinna sitter vid ett bord, kvinnan håller upp händerna i fredssymbolen.
En man och en kvinna sitter ner.
Fyra små barn klär sig i svart och röd bröllopsklädsel spela på golvet.
En person på en cykel drar en vagn full av pinnar.
En man i en färgstark skjorta klädd som en clown.
En liten flicka i klänning sitter på trappan för att äta mellanmål.
Kvinnan som bär en fluga går längs New Yorks gator.
En grupp gatutrummisar spelar medan några åskådare dansar.
En man i halmhatt som bär ryggsäck rider på en motoriserad skateboard.
Tre damer låg på en strand som vetter mot havet.
En person lyssnar på musik över sina hörlurar medan han går nerför en övergiven gata.
En kille på ett kontor lagar kaffebryggaren.
En man i röd tee-shirt styr sitt cykelliknande fordon på en gata i Santo Domingo.
Två kvinnor går nerför en trottoar.
En ung dam i ljusblå kläder som går längs en vackert designad trottoar.
En kvinna i solbränna går nerför en livlig trottoar.
Två poliser ser män på en motorcykel, med en vit is bröstet på den också, bär hattar
Mannen sitter i gul bil i solen, torka pannan.
En man tittar bakom den skyddande buren på ett tungt maskineri medan han bär skyddande hörlurar på huvudet.
En man och en kvinna som sitter, med en man som står till vänster.
En kvinna i grön topp och orange shorts går på gatan.
En man knuffar sin blåmålade snacksvagn genom gatan.
En kvinna och 2 små barn leker i sprinklers från marken.
Folk tävlar för att fånga tunnelbanan i skymningen.
Män och kvinnor vid bord med drinkar på akterdäck på en båt förtöjd i en marina.
En man stirrar ut över en bangård.
Fyra personer står bredvid några cyklar medan en av dem poäng.
En man på scenen framför en flagga som talar in i en mikrofon till en publik.
Tre personer står på en matta och en har en sele på.
Män går nerför en gata och spelar trummor.
En kvinnlig anställd på en fiskmarknad väger en vara på skalan.
En man köper sina grönsaker på marknaden.
Två bruna hundar leker tillsammans i vattnet.
Män som promenerar i ett tegelmålat, ljust upplyst affärsdistrikt.
En man och kvinna som är intima i ett stort tomt rum.
Två barn på en båt tittar av, blå våningen.
Ett litet barn som ler och tittar utanför fönstret.
En skara människor tittar på något utanför en Gap-butik.
En äldre kvinna får pengar från plånboken i en annan kvinnas monter på gatan.
En man i khakibyxor och en kvinna i kjol korsar en gata.
En ung flicka i kamouflagefärg håller i en rosa skylt.
Två kvinnor i mitten av gatan pratar.
Två kvinnor i kjolar står tillsammans bakom ett metallstängsel på en allmän gata.
Två personer står och pratar med varandra.
Ung asiatisk pojke sätter sig ner och läser en bok på en bokmässa när en kvinna tittar på.
En kvinna tittar på sin mobil medan en man tittar på henne.
En flicka i vit skjorta, som går bredvid sin cykel.
En grupp människor sitter framför en lägereld.
En kvinna med sneakers och en kjol sveper ut en lagerbyggnad.
En grupp människor marscherar i en parad som viftar med flaggor.
En kvartett ungdomar, kanske spanska eller portugisiska, bär röda bandannor, medan en iögonfallande inte gör det, promenerar nerför en boulevard.
Det verkar som om de förbereder sig för mötet.
En grupp ungdomar sitter i baren och umgås.
En humvee visas mitt på ett torg.
Två kvinnor sitter i gröna stolar och en liten pojke i röd skjorta kastar ett tecken.
En man i blå Speedos håller i svarta glasögon.
En grupp människor i vita skjortor och röda bandannor samlas tillsammans.
En massa människor tittar på en anslagstavla på kinesiska.
En ung man i kostym sitter på en buss med huvudet nere.
Ett litet barn som bär en gul skjorta står på trottoaren.
Flera personer tvättar sig själva med hjälp av duschar på stranden.
Grupp med gula och orange skjortor ridande mountain bikes.
En man med glasögon och en ung flicka som ler mot kameran ger flickan ett fredstecken.
Tre tjejer rider på en berg-och dalbana.
En liten pojke i grön skjorta äter chokladglass.
En man i grå t-shirt sitter mot ett trottoarträd.
En liten flicka med svarta grissvansar rider en rosa cykel med träningshjul.
En liten flicka som bär en vit blus står efter böcker.
En man i blå jeans som sitter framför en affär.
En kajakpaddlare går genom några kurviga forsar.
Mannen är i en gul kajak i grova vatten.
En man står över en bås med en stol täckt av en sporttröja.
En kvinna sjunger på scenen när en man spelar ett instrument i harmoni med sin sång.
En man i blå rock spelar gitarr under ett träd.
En grupp äldre människor som besöker en marknadsplats nära en tupp.
En kvinna väntar på ett tunnelbanetåg.
Två små pojkar med skedar som rör om i två metallpannor.
Man drar en vagn full av hinkar, moppar och kvastar.
En kvinna med starkt rött läppstift, solglasögon och en röd rutig skjorta tittar mot kameran.
En man bär röd skjorta och väst.
Kvinnan i Jacket med huva upp promenader ensam på trånga gatan.
Två kvinnor i klänningar som går längs trottoaren.
En kvinna vid ett utomhusevenemang har en broschyr i handen.
Band på scenen och folk som tittar på skärmen.
En skara människor tillsammans i ett område.
En kvinna med rullande bagage väntar på en trottoar.
En gammal man med blå skjorta står mot en vägg.
En man på ett kontor leker med ett barn
En man i orange overall använder en rulle för att täcka graffiti.
Mannen i grå skjorta och svarta byxor står framför en butiksfront.
Tre parkerade taxibilar med två parkerade polisbilar bakom sig.
En man i en läskig potatissäcksmask.
En kvinna tar en paus från att sopa upp en trasig gryta för att titta ut genom fönstret.
Äldre män koncentrerar sig medan de spelar en omgång Dominoes.
En man och en kvinna ligger tillsammans på en gräsbevuxen parkfält nära en strand.
Folk går förbi Starbucks Coffee store med gröna markiser.
En man och en kvinna som håller hand när de går.
En man på en cykel leder en häst och ryttare i ett landsbygdsområde.
En butik med två män utanför, en man in i butiken, och motorcyklar synliga på höger sida av ramen.
En man i en fluga arbetar med trä.
En man i svart hatt pratar med en kvinna med en djurskjorta.
Flera grupper av fotgängare på en stad gata under dagen.
En kvinna i en grön jacka står vid en vägg full av konstverk, framför en butik som visar kläder och skor.
En kvinna i en blå jacka som går ut.
En man som spelar fiol står framför en annan man som spelar dragspel.
Två män i halmhattar står vid en höhög på en livlig gata.
En man i skinnjacka sitter på ett staket vid stranden.
Kvinna i klackar och kjol tittar på produkter.
Blond kvinna i blå outfit hänger på golv kudde vid utsidan bord ensam.
Pojke som leker i vatten kommer från fontänen.
En flicka som bär rosa går förbi en väggmålning av en flicka med rosa hår.
En man i svart skjorta som sitter vid ett restaurangbord och sms:ar.
Två kvinnor i vita klänningar poserar på en filt för fotografier mitt i en park.
Folk samlas på ett gathörn i sommarkläder.
En man med latexhandske och svart skit står framför en Chevy van.
Två kvinnor bredvid en scen av människor spelar instrument
Folk går och en dam tittar på hennes mobiltelefon medan de går i en stor stad och handlar.
En person ligger på en blå filt på en trottoar.
En man och en kvinna kommer nerför en rulltrappa.
En kvinna med långt hår som sitter på en betongbänk.
En kvinna bär ett barn, bär gröna hörlurar, på ryggen
En smet förbereder sig för en swing under en omgång cricket.
En person som sitter framför en laptop och många elektriska delar.
En man som fiskar vid en liten brygga vid solnedgången.
Ett flygplan står med en gotisk byggnad på baksidan.
En liten unge som leker i vatten.
En man med solbränd jacka går förbi en kvinna i hästsvans.
En man som står framför en glasdörr.
En grupp människor samlas i en protest mot våldet i Mellanöstern.
En asiatisk kvinna som hade ryggsäck och flinade över axeln.
En kille i khakis och sandaler är på en tvättmatta.
En man knuffar ner många kartonger med bröd på gatan.
Ett flygplan som flyger över ett staket med några åskådare som tittar på det när det närmar sig sin landning.
En ung pojke som övar på att slå en baseball från en tee.
En man och en kvinna som går uppför en gräsbevuxen slottsfil.
Folk väntar på ett tåg vid tunnelbanan.
En grupp människor står på trottoaren framför flera butiksytor, med en vagn parkerad nära dem.
En äldre man spelar fiol på gatan.
Människor passerar tiden i en stad i ett mellanösterländskt land.
Man i vit skjorta står på gatan med säljare och massor av människor.
Ett plan flyger lågt över ett gräsområde där en flicka sitter i en fällbar stol.
En man som bär svart sitter utanför under palmer nära gröna och blå stolar.
Tre unga flickor står utanför nära ett staket leende mot kameran.
En grupp människor i vita uniformer bygger mänskliga stege.
En man pratar på sin telefon bredvid vit tegelvägg med blå färg stänkt på delar.
Ett blond barn gömmer sig bakom en trästolpe.
En ung dam läser en bok medan hon sitter ute vid foten av en palm.
En blond kvinna poserar med två personer målade för att se ut som statyer.
En del människor sitter, en del står på en trottoar.
En man i kostym röker och pratar i telefon.
En blond kvinna i en tank topp och shorts sätter sin fot i en fontän.
En man sjunger och flickan spelar ett instrument.
En bild av duvor som lyfter med en ung flicka i den avlägsna bakgrunden.
En person som håller i en platt låda står nära två personer som sitter ner.
En manlig simmare i en blå Speedo baddräkt anpassar sina glasögon.
En man i en tanktopp tittar på en kvinna nära en vattenskulptur.
Två äldre kvinnor sitter på en bänk och samtalar.
Två unga pojkar vandrar genom en folkmassa med ljusgula skjortor.
En man med hatt, vit skjorta, byxor och skor sover på en parkbänk.
En man som väntar i tunnelbanan bredvid bussen och läser tidningen.
Ett barn som springer genom vatten utanför en park.
Två kvinnor och två män som står under ett regntäckt tält.
Den här unga flickan bär en röd och svart rutig skjorta.
Grön cykel sitter utanför på trottoaren på displayen.
En man som står på en scen och spelar gitarr och en munspel som vinkar till publiken.
Flera asiater framför butikskoncept.
En man i blå skjorta sitter på en dörr och pratar på sin mobil.
En liten pojke och hans far säljer snökoner från deras spårvagn.
En flicka läser och lyssnar på musik på en buss.
En välklädd kvinna handlar framför en affär.
En fullsatt stadsgata med fokus på en äldre man som spelar gitarr.
En man slumrar till ovanför några gröna glas.
En person i shorts med en tatuerad kalv håller kopplet på en stor vit hund i en blå väst.
En man avfyras i luften från en flotte.
De sex människorna är i en blå flotte i vattnet och en person flög ut ur flotten.
En man i en ärmlös skjorta som vilar vid trottoaren.
En liten flicka och pojke på baksidan av en cykel väntar på pappa att trampa.
Två svarta män står framför en ljus stolpe.
Tre personer kantade på gatan och skuggade sig själva från solen med paraplyer.
En man vill köpa flaskor på en marknad.
Folk tittar på en man som klättrar på ett rockansikte.
En kvinna som bär en Wonder Woman-dräkt och en röd jacka.
En äldre kvinna som bär hatt och rosa skjorta njuter av en cigarett.
En man som bär på en jättelik bananleksak går på gatumässa med ett litet barn som håller hans hand.
Mannen tittar ut ur sin blå bil och håller ut en trasa genom fönstret.
En grupp människor ro på en sjö.
En gammal kvinna med vit skjorta och gröna shorts står på en trottoar.
En man i vit t-shirt tittar bort från kameran.
En grupp på fyra män som diskar och torkar i ett kommersiellt kök.
Två manliga studenter städar i ett labb med stolarna uppvända på borden.
En pojke bär rosa slips och en annan pojke bär en flickas klänning, och många människor i bakgrunden.
En man i svart jacka och hjälm vid handen poserar med ett leende.
En ung pojke i cowboyhatt och en blå jeansjacka som sitter i en barnvagn.
En svart kvinna i randig klänning som sitter på en blå bänk.
En person står bredvid ett träd med solen skiner genom löven.
En pojke och hans far går i cowboykläder.
En man i svart skjorta springer nerför en livlig trottoar
En äldre herre som talar på ett podi.
Två unga pojkar med shorts leker utomhus medan en polis vaktar.
En gammal man med glasögon framför ett podi.
Ett barn i röda byxor som håller en metallkorg bredvid ett annat barn i en blå jacka.
Två damer visar tillgivenhet som leder till en kyss.
Det finns en grupp av många vuxna runt en falsk pirat fartyg klädd som pirater.
Gammal person som går längs trottoaren bredvid en vit byggnad.
En röd vintage bilparkering framför Karlova 25.
En tonårspojke som bär mössa ser irriterad ut
En leende medelålders man som bär överstora röda solglasögon och en färgglad mönstrad skjorta sitter i gräset framför en blågrön bakgrund.
En liten röd och vit tävlingsbil tävlar under loppet.
En man som bär keps och glasögon håller på att fästa sätet på en cykel.
En kock lagar mat på en wok på en utegrill.
Ett mans- och kvinnopar går förbi väggen målat med figurer av människor och graffiti.
En person sitter på en klippavsats med utsikt över en vattenförekomst.
Ett grönt föremål med ljus hängs upp över en trottoar där tre personer går.
En man håller sitt tal.
En man med en vandringsutrustning knyter sin sko i skogen.
Flera kvinnor utför en dans på ett formellt evenemang.
En asiatisk kvinna på en fullsatt plats som gör sig redo att knäppa en bild
En grupp barn går i sanden.
En kvinna som torkar pannan av en annan kvinna, sitter ner bland en skara av kvinnor, dricker från en flaska.
En man med glasögon som spelar en silvergitarr.
Tre vandrare står nära och på en träkonstruktion som delvis består av stockar.
En bar med en man och en kvinna som pratar
En man i gräddskjorta sitter på en utomhusrestaurang med en svart bil bakom sig.
En man med en stor mohawk och DIO skjorta manipulerar en mobiltelefon.
Brun, svart och vit hund som står på en sandig sluttning.
En grupp människor i gröna skjortor som går längs en vacker strand.
En man i kostym skakar hand medan två andra herrar tittar.
Fem personer poserar för ett familjefoto.
En kvinna som håller i ett rött parasoll tar en bild när hon tittar över en vägg.
En kvinna och en man som bär en rosa kylare.
En pojke i en blå tanktopp spelar basgitarr med en fot i luften.
Två personer på en vit strand, en har en mycket lång pinne.
En ung flicka i baddräkt som dricker ur en grön glasflaska
En kvinna som bär shorts och sandaler korsar gatan med gula taxibilar i bakgrunden.
En grupp människor som går utanför en nöjespark mitt på dagen.
En skara människor som står utanför en byggnad.
En ung man som bär en röd t-shirt och svarta byxor utför en framhjulsställning på en cykel.
En turist går under skuggan av en byggnad.
En kvinna i en lila halv skjorta och en kjol som går nerför en gata.
Människor utanför på ett fält skördar något.
En ung man i randig skjorta håller upp en stock i en park.
Fyra barn leker i en swing set.
En äldre asiatisk man som tittar ut ur en byggnad med solljus på väg in.
Två män i solglasögon går nerför gatan.
Två kvinnor med alkoholhaltiga drycker i sina händer samtalar med varandra.
En man som sitter ner och läser en bok.
Glasfönster visar upp en modell av en man som sitter och bär svart.
Damen tar bilder på statyn.
En man i vit skjorta och svarta byxor står vid sidan eller vägen.
Ett ungt par med barnaffärer på en liten smörgås och kafé.
En man med mustasch och gitarr sjunger för dricks på gatan.
En person står under en stadsljusstolpe på en trottoar på natten.
En blond tjej som har ett samtal med sin brunettvän på en utomhuskonsert i regnet.
En grupp människor tänder lyktor.
Grupp av män och kvinnor som sitter på lådor och hinkar i ett utrymme med medel ljus och mat.
Två bilar och tre män står bredvid en lastkaj.
En kvinna i ett förkläde rengör ett bord som är omgivet av olika färgade stolar.
En man med långt hår lutar sig mot en kedja samtidigt som han håller en bild.
En man står inne i en dörröppning som är i en vägg målad med en väggmålning av en kvinna.
Tre personer tittar på en fjärde rita en krita porträtt på gatan.
En grupp människor samlas utanför runt en staty.
En kvinna som sätter smycken i fönsterfönstret.
En man cyklar genom en smal väg mot ett torg som gränsar till ett slott med ett blocktorn.
Två personer går över en stig mellan byggnader.
Ett par går under en båge på en smal gata med balkonger.
En ung pojke sitter ute och säljer för pengar medan han spelar dragspel.
En kvinna går nerför gatan med hörlurar i öronen bredvid en man i kostym.
En svart tröja som bär en lila väska på gatan.
Två kvinnor sitter och tittar åt samma håll.
En afrikansk amerikansk dam som har en korg på huvudet.
Detta foto innehåller en staty av en man och en kvinna som går med en blå skjorta som går bakom den.
Flera personer promenerar genom en park med många träd.
En kvinna på en gata tar ett foto medan folk går förbi.
En man lagar något på spisen.
1 man står och flera människor sitter och väntar på ett tunnelbanetåg.
En manlig konstnär som ritar med krita på gatan.
En upptagen pizzabutik ligger på ett mycket trafikerat gathörn.
En polis kör sin motorcykel längre ner på gatan.
En grupp orientaliska ungdomar står utanför dörren till en affär.
Detta är en bra karta för turister.
Två kvinnor på tunnelbanan helt hänförda med sina prylar.
En man går förbi ett graffitierat område.
En grupp på tre kvinnor och en man tittar in i ett skyltfönster.
En man i en läkarrock kommer från en byggnad.
En man och ett barn är tillsammans med ett blått nät framför dem.
En kvinna som handlar frukt på en utomhusmarknad.
En man som säljer glass från en vagn till ett litet barn på gatan.
En lantbrukare i utbildning pekar över barriären vid en boskapsauktion.
En dam med glasögon som spelar saxofon framför en affär.
Fyra tjejer sitter i en bubbelpool.
En man står på en transportplattform med hörlurar och en handhållen elektronisk apparat.
En man i gul skjorta läser en bok.
Man med randig ryggsäck rullskridskor nerför en upptagen aveny med andra rullskridskor.
En man sitter på en fyrkantig sten och äter sin lunch.
En asiatisk skolflicka i en typisk skolflicka uniform, mörk pullover, rutig kjol och knästrumpor med öre loafers.
En kvinna i en röd halsduk som går genom en ingång på en gata.
En flicka leker med leksaker i ett badkar med vatten.
Två personer lagar mat på en solig dag för andra.
Medan mannen väntar på ett tåg läser han en bok.
En afrikansk amerikansk kvinna plockar tomater i en trädgård.
En medelålders man med glasögon och en medelålders kvinna ser både grinig och upprörd ut.
En spansk gitarrpolare och en damdansör som uppträder på scenen.
En liten flicka gör ett handstöd på en studsmatta
Ett litet barn med turkosa shorts som står nära ett stort träd.
En grupp kvinnor alla på liknande sätt klädda marscherar med ett stort föremål på sin högra sida.
En publik som njuter av en konsert.
En skara människor samlas runt Oxford Circus Station i London.
Folk sitter och ser på när en gatuartist sjunger.
En ung man som bär en grön skjorta tar hand om en tomatplanta.
En man i grön skjorta med en boxskärare omgiven av grönsaksväxter.
En kvinna som bär glasögon sitter vid ett bord med glasögon, en flaska och en fågel på.
En man och två barn tittar på en kamera.
En ung kvinna går nerför gatan förbi ett fönster som är täckt av tidningen.
En bronshudad kvinna går en gångstig i en form som passar klänningen.
Två äldre män sitter på skotrar framför ett Koffee Cafe.
Tre personer sitter på trottoaren på vägen.
Många människor och bilar går förbi ett kafé i hörnet av gatan.
En grupp duvor går på en trottoar.
Tre personer försöker öppna en stor dörr till en stängd butik.
En hektisk dag på stadens gator.
En äldre kvinna sitter vid ett restaurangbord under en skylt på väggen och läser "Oh boy mammas pannkakor!"
Fyra personer går nerför en trottoar - tre mot kameran en bort.
En ung man som jobbar hårt och sopar golvet.
En kvinna sprang förbi ett par människor som satt ner för lunch.
En man i uniform korsar en gata.
En kvinna går förbi en gammal bagelbutik.
En mor och ett barn som går i regnet i ett grönt område.
Äldre fiskare roddar en grön båt som står upp för en lugn flod.
Tre segelbåtar går nerför vattenvägen i ett tropiskt slätt vattenområde.
Byggutrustning och arbetstagare i en stad utanför USA
Det finns en äldre kvinna med en ljusgul skjorta som står på en trottoar och tittar in i en affär.
En man drar sitt matstånd tvärs över gatan.
En kvinna dansar i en färgglad klänning, engagerad i en vresig dans som hennes äldste lärde henne.
Två flickor med klänningar står på en murad trottoar.
En man i en folkmassa framträder i en stadsscen med en mestadels svart dräkt med en grafisk bild på sin skjorta.
En man drar på ett rep i landet.
En kvinna går på trottoaren med en annan person som följer efter henne.
En omtänksam kvinna går nerför en storstadsgata.
En man sätter sig ner för att vila på en fullsatt gata.
Barn kvinna och man i en park tittar runt i en park
En äldre man hugger ved bredvid ett stort träd på en åker.
Personen i vit T-shirt går.
Kvinnor med falskt blod och smink över hela ansiktet, bröstet och halsen.
En man steker gladeligen kinesisk mat.
En gatumusiker i blått, med en cigarett i munnen och en stor gitarr i händerna.
En gata med gatubelysning och busshållplats.
En grupp buskiga håriga människor går nerför en regnig trottoar.
Kvinnor i rosa klänning med vita prickar stående på sten bas shoo-shes de i utsikt.
En kvinna med en crossbody svart handväska går nära en trappa med silverräcke.
Två solbadande människor sitter på en bänk framför en brud och brudgum.
Ett litet barn i orange klänning tittar på graffiti av en afrikansk amerikansk baby.
En Toddler med en blå designskjorta och grå kort valsning med sin familj.
En man med grå kula går bredvid en rödhårig kvinna i en långärmad blå jeansskjorta.
En röd metallskulptur omges av ett stort antal människor.
Två kvinnor vid stängslet medan ett barn springer mot dem.
En vacker ung kvinna håller i sin handväska.
En kvinna i svart skjorta skapar konst på trottoaren.
En söt liten unge med lite grönt klistermärke på näsan.
Tre män i vita skjortor poserar för en bild utanför en lokal butik.
En kvinna i jeans shorts poserar för fotot.
En man som bär solglasögon ses på en solig dag bredvid en skulptur i en park.
En man med en vit hjälm i publiken.
En kvinna som står i ett rum som är vitt med siffror i en cirkel runt henne.
En man står på stranden.
En grupp judar viftar med flaggor för att fira sin religion.
En naken man inlindad i ett nät som ligger på några klippor på havssidan.
Röda kinesiska lyktor och banderoller på kinesiska hänger en livlig gatuscen.
Vi kan se blod på baksidan av den här mannen
Folk bläddrar igenom objekt på en öppen marknad.
En del kaukasier tycks tillaga mat och dryck.
Solglasögon sitter på ett bord med familj på en brygga i bakgrunden.
En kvinna som står framför en affär som heter La Perla.
En grupp människor samlas utanför medan en man i svart skjorta och glasögon går mot kameran.
En grupp slumpmässiga fotgängare tittar på något utanför kamerans räckvidd.
En person springer på en skogsgata med solen i bakgrunden.
Den skäggige mannen i hatten höll kameran i båda händerna och väntade på nästa skott.
En välklädd äldre kvinna som står framför en buss dekorerad med bilder av lila blommor.
Nån i blå jeans och en blå luva som täcker ansiktet och fixar en cykel.
En man i en ljusrosa polotröja håller en flagga utspelad i luften bakom honom.
Folk på en karneval deltar i en skjuttävling.
En man med smink i ansikte och hals som ser ut som blod och sår.
En äldre man ser en yngre man grilla olika maträtter.
Ett par försöker hitta den plats de vill åka till.
En man sitter och skriver vid ett bord som är uppställt på en trottoar.
Tre män står medan en annan står bredvid dem med en tidning.
Smickrande brunett med rödhårig klänning deltar i en parad.
En spansk kvinna i ljusa färger klädd för en parad.
En tatueringskonstnär som gör en kvinnotatuering av en ros
En man och en kvinna står på en båt medan mannen fotograferar.
En kille med vit skjorta tar en bild.
En vacker kvinna i persikoklänning går nerför en tegelgata på natten.
En svart streetdansare uppträder för en massa människor.
Ung pojke sparkar en röd och vit fotboll på en gräsbevuxen åker
En man som får magen tatuerad av en tatueringskonstnär.
En man och en kisande kvinna tittar på något på en skärm.
En kvinna i en violett skjorta står vänd mot en ung man.
En man i vit skjorta och khakibyxor kollar sin mobil framför ingången till en byggnad.
En tatueringskonstnär som jobbar på en tatuering.
En tatueringskonstnär som gör en tatuering på en underarm.
En man i jeans får en ny tatuering.
Två unga pojkar spelar några instrument vid vattnet.
Ett suddigt foto av ett par på en bänk som ser andra människor spela.
En kvinna ser en dinosaurieskulptur i metall genom ett blått teleskop under en molnig dag.
Äldre kvinna som försöker blockera solen med handen.
En man och en kvinna klädd i svart är rullskridskor.
Två unga kvinnor går och pratar.
Kvinnor i färgglada klänningar dansar nerför gatan under en parad.
En frisbee kastar en skugga på hunden.
Konstverk av ett litet barn och hans hund har utsikt över en lugn trottoar och en man som sover mot sidan av en byggnad.
Två personer klädda i superhjältedräkter står på stans gata.
En kvinna som står bredvid en fotograf ger ett papper till en man i grön skjorta.
En tjej åker rullskridskor längs en gata medan hon pratar på en mobiltelefon.
En ung pojke står på en idrottsplats och håller i en sportutrustning.
Två unga damer går längs gatan tillsammans.
En kvinnlig trafikofficer som leder trafiken i en livlig stadskorsning.
Gentleman står på en trottoar och tittar på en byggnad.
Det här måste vara en av de bästa restaurangerna på östra sidan!
Pojke i röd skjorta med kamera.
En man går på gatan när han börjar passera glasfönstret i ett företag.
En stav besättning, av fem, reparerar en väg.
Här är en bild på en kvinna som ler mot kameran och röker cigaretter vid en middag med levande ljus.
En man som spelar gitarr medan en kvinna kollar ugnen.
Två kvinnor står vid en stor serie av skyltar som säger "Le Cafe Marley" i en hall med ett mycket högt och utsmyckat tak.
Tre kvinnor går nerför en trottoar nära en bistro.
Två män spelar schack i parken medan två andra ivrigt väntar på sin chans
Folk går längs en gångväg omgiven av byggnader.
Ung man ser på som en annan man som sitter på ett staket lindar sina ben runt en hona i en zebra stil tank topp och kjol.
Tjej i kort svart klänning Blåsa en gigantisk bubbla för en publik utomhus.
En kvinna och barn sitter på trottoaren vid ett träd medan en kille lurar runt i bakgrunden.
En man i svart huk med folk som går tvärs över gatorna.
En man i vit skjorta pratar med en kvinna i grön blus på gatan.
En man som håller i ett ljus med huvudet lutat mot en staty.
En kvinna i solbränd topp och jeans sitter på en bänk med hörlurar.
En man och en kvinna som går nerför gatan med en shoppingväska.
En grupp människor sitter på en vägg ovanför en stor basrelief-skulptur och reflekterande damm.
Två vackra flickor visar sina praktfulla kroppar.
En man i hatt står vid ett hörn framför en rad cyklar.
Kvinnor njuter av drycker på en restaurang utanför.
En kvinna poserar ovanpå en skoter medan en fotograf förbereder sin kamera.
En ung kvinna tar bilder medan en folkmassa salonger på en grön gräsmatta.
En kvinna med blont hår och svarta byxor övar sina karaterörelser i en naturskön park.
En man står framför ett väl upplyst fruktstånd.
En person som bär solglasögon och en ljus orange skjorta går nerför en våt trottoar.
En man och barn sätter upp en monter för att sälja smycken.
En gammal byggnad med en lång hall och glastak.
Två poliser på skridskor står nära en annan man.
En man i hatt och en pojke i hatt sitter utanför Louvren.
Två män tar bilder med sina kameror utomhus.
Folk njuter av det svala vattnet från fontänen på en varm dag.
Två män sitter på kanten av en vattenpöl.
En man klädd i alla vita kläder står framför en grå vägg, armarna korsade.
Unga kvinnor och män klädda i kostymer sittande och stående.
En bergsvandrare gräver biffar i snön.
Folk sitter på en buss.
En man sopar vägen framför en vägg med graffiti och två lägenheter mot den.
HO King producerar en butik som erbjuder snöärter, broccoli och napa.
En äldre asiatisk man väntar på att någon skall ge honom service vid en matdisk.
En man visar upp olika typer av skaldjur på en pinne, däribland sjöstjärnor.
Två män undersöker ett cykeldäck medan en kvinna i bakgrunden lutar sig mot en vägg bredvid en gryta med pelargoner.
En man som sitter på en bänk bredvid sin cykel.
En grupp människor som står nära en båt på en vattenförekomst.
En kvinna i klänning pratar i telefon.
En dam sitter på slutet av en pir högt ovanför vattnet.
Två kvinnor pratar med en man i en keps.
Tre vuxna står framför en skylt som säger "rösta" och en amerikansk flagga.
Bagagevagnarna är uppradade och redo att flyttas.
En kvinna står i ett bås, bär och orange väst, erbjuder ett kreditkort och ler.
En kvinna går hundar på en väg som ligger i staden.
En kvinna lägger sig på en flytande plattform mitt i en vattenförekomst.
Två unga vuxna utanför, med många träd i bakgrunden.
Två stora kukar syns utanför restaurangen el pub restaurant.com.
Två män går sin kanot genom skogen.
En man i en kanot sitter på en lugn sjö omgiven av grönskande lövverk.
En man och en kvinna som visar ett litet barn hur man använder ett vapen.
En man som spelar en unik fiol medan han tittar upp i taket.
En violist som spelar bredvid en reklamskylt
En man i vit skjorta och långt hår som spelar elviolin.
En violinist som spelar musik i tunnelbanan i New York.
En person bär sin vita kanot nerför en stenig stig medan en svart hund i en röd krage klockor.
Mannen som bär allt svart sover på sin röda motorcykel.
Ett litet barn med en hatt på att leka med en bubbelmaskin.
En präst med buskigt skägg som äter snabbmat.
En man som bär en blå och svart rutig överskjorta säljer ekologisk frukt till en man i en grå poloskjorta.
En kille som spelar dragspel med hatt på.
Jimi Hendrix har blå kläder när han spelar gitarr.
Det finns två bruna hundar som leker ute på fältet.
Publiken tittar på hästen, stirrar på cowboyen när han lämnar arenan och undrar vad som kommer att hända härnäst.
En kvinna som går på en förortsgata.
En man undervisar små barn om att laga cyklar i en park.
Musiker uppträder utomhus för pengar.
Gatorna i en Chinatown ser likadana ut är upplysta med ljusa färger.
Några grupper går nerför trapporna.
Det finns flera personer som antingen sitter på bänkar eller går genom vad som verkar vara en tegelväg med träd som kommer upp från olika cirkulära öppningar i vägen.
Flera asiatiska fotgängare går runt en silvertaxi van.
En liten flicka i en röd print sundress gick genom en utomhus konstnärsutställning.
Ett fotbollslag ses göra pjäser, blockera, fånga och springa.
En man tittar på en karta medan en kvinna i solglasögon tittar upp.
En man i vit skjorta läser en karta.
En afroamerikansk man i grön skjorta och solbränd jacka.
En man i lila skjorta och blå jeans spelar munspel av en röd buss.
En grupp män, kvinnor och ett barn går i en grupp.
En kvinna kramar en man.
En dam i vitt sitter på en matta med en boll i handen.
En asiatisk marknadsplats är öppen för affärer på natten.
En kvinna tittar på medan en annan kvinna tar en tallrik mat.
Två män och en kvinna i ett band som spelar en låt.
En ung flicka och en pojke simmar under vattnet i en pool.
En hund i en bil.
En grupp människor passerar en tunnelbanestation.
En blondhårig mor håller sitt nyfödda barn.
Ett litet barn får bad i ett plastbad av en vuxen som bär gummihandskar.
Kvinnorna tvättar det nyfödda barnet.
En topless kvinna vaggar sitt nyfödda barn svept mot bröstet på sjukhuset.
En skara människor går genom en livlig gata.
Äldre kvinna i en ljus lila skjorta, sitter i en stol, håller ett barn.
En man och två unga pojkar sitter på en sten.
En liten pojke och en liten flicka som leker i en fontän.
En upptagen kvinnor i svart och vit färg klänning korsar vägen.
En mamma och dotter går uppför trappan när en kvinna bär en huvudduk i närheten av en soptunna.
En fransk cykelhytt utan passagerare som sitter vid en trottoar.
En ung flicka skrattar och jagar duvor på gatan där andra människor går i närheten.
En turist tar ett foto av något högt.
En kvinna håller en mycket stor mobiltelefon upp till örat.
En man och en kvinna, båda klädda i solglasögon, tittar upp mot himlen.
En man med en shoppingväska och en kvinna tittar på en kamera.
En kvinna som håller i en svart plastpåse håller en digital kamera ovanför.
Ung man som sitter på fäktning framför vackra blommor trädgård håller två unga damer på knä.
En dam går uppför trappan från tunnelbanan.
En utsikt över en skara människor som går längs sidan av en flod.
En väl upplyst reklammonter visar upp olika filmaffischer.
Två olika grupper av människor samtalar framför Shakespeare och Company butiken.
En man kör en vit skåpbil sprejad med graffiti.
En man med ett protesben sover framför ett lager.
En person ligger i en sjukhussäng.
Antingen gör sig en dam redo att gå till eller så har hon precis slutat opereras och födas.
En medelålders kvinna håller i ett barn.
En nyfödd är insvept i en randig filt medan någon rör vid den med båda händerna.
Man håller gråtande bebis i stolen nära fönstret.
En läkare och hennes patient ler klart som ett spädbarn sjuksköterskor vid patientens bröst.
En man i svart skjorta håller ett barn.
Två män sitter där ute och tittar på en tidningsbild av en kvinna i bikini.
En äldre herr med mörka byxor och en vit skjorta går genom en park.
En stadsgata med några förbipasserande, med en stenblocksvägg med graffiti på.
Åskådarna fascineras av en man som jonglerar med flammande stavar medan han rider en enhjuling.
En man står utanför en vacker byggnad med neongrön byggjacka.
En dirigent ger ett barn en rundtur i tåget.
En man är på en avslappnad cykeltur under dagen in till stan.
En kvinna med solglasögon sitter under ett rött paraply
En flicka med lila klänning och en flicka med röd klänning springer runt utanför och ler.
Flera grupper av människor går i en vacker park.
Telefonkiosker upptagna av några personer.
Två blondiner delar ut flygblad och ballonger på en livlig gångväg.
En man på en BMX cykel utför ett trick på ett hopp.
En taxi i en korsning i centrum.
En polis i Madrid i Spanien stannar för att tala med en äldre kvinna.
En motorcyklist rider förbi ett asiatiskt snabbköp.
En kvinna med parasoll rider sin rosa cykel nerför gatan.
En familj på tre personer tittar på när män i kostym passerar förbi.
Två personer i blå skjortor tar ett foto av sig själva som en kvinna i en halsduk passerar dem.
Ett par promenader längs en trottoar.
En man med långt vågigt hår spelar för violin.
Två män på en gata, en med röd flagga.
En grupp ungdomar står framför och rör vid en svart, rostig metallstruktur.
En man i hjälm hänger på sidan av ett transitfordon.
En skallig man tittar ut över en skara människor.
En grupp människor samlades runt en monter och sålde öl.
En grupp människor går framför en stor stenbyggnad.
Människan samlar papper nära en struktur av trä täckt med papper och graffiti.
En person i lila klänning, svart hatt och rosa halsduk kör på en väg.
En man i shorts och en orange skjorta sitter på bakluckan på en lastbil och undersöker en telefon.
En man sitter på ett tåg och lyssnar på musik.
Två unga flickor går längs en gångväg med ett paraply.
En person med svarta handskar och vit hatt står och justerar sin halsduk.
En ung man går lättvindigt nerför gatan framför några träd.
Två kvinnor med långt hår och hästsvans joggar längs vägkanten.
Ett gäng seniorer samlades i ett område.
En person i en cowboyhatt rider på en solbränd häst.
Två personer som sitter på en parkbänk och tar en tupplur.
En tjej med blont hår är kopplad till band av många färger och njuter av någon form av firande.
En man med svart ryggsäck knäböjer över en hög med affischer.
En stor skara människor väntar framför en stor talare.
En rad lastbilar går nerför en mycket trång gata.
Folk som bär mönstrade t-shirts firar några festivaler med färgglada ögonkläder
En skäggig man balanserar en silverboll på ena handen.
En liten unge i svart som leker i en fontän.
En ung man som bär ryggsäck bär en vit kartong.
Tre personer av asiatisk härkomst står i en halvcirkel och pratar medan en tjej sms:ar.
Folk går på en fullsatt gata.
En kvinna i klänning och cowboystövlar går bredvid en annan kvinna i en svart t-shirt.
En kvinna i lång kjol och en man går nerför gatan.
En grupp män uppträder på trottoaren med sina gitarrer.
Två unga flickor poserar för en bild bredvid vattnet.
Två skjortlösa små pojkar, den ena lutar sig mot den andra, står på en stor sten framför några träd.
Strandpromenaden är mycket ljust upplyst av restaurangskyltar på natten.
Det ena barnet tar bort munstycket från det andra som får honom att gråta.
En kvinna bär påfågeldräkt.
En solig dag sitter en man på stenar och röker bredvid en vattenförekomst.
En man i blå jacka cyklar på trottoaren.
En grupp elever är utanför, väntar, framför en gul skolbuss.
En kvinna som tittar på sin telefon och håller i sin pomeran.
Två kvinnor väntar på trottoaren framför en stor reklambanner.
Fyra personer står utanför en närbutik.
En rödhårig kvinna sitter på en bänk i randig kjol och bruna skor.
En man njuter av en smörgås från Subway.
En man som går ifrån en rulltrappa medan en kvinna kommer upp för rulltrappan.
En pojke står i en båt, håller upp en fisk till kameran och ler.
Ett countryband på scen som spelar musik i gult och rött ljus.
Sex personer på nån sorts konferens.
En man med vit skjorta, bruna skor och blå strumpor läser nära andra människor och högar av böcker.
Asiatisk man i vit tank topp äter av en stor asiatisk politisk gobeläng.
Den lilla flickan såg med vördnad på synen.
Gatuvy över Orient Hotel.
En man på en röd cykel som släpar en vagn bakom den.
Folk går på Times Square i New York.
Två hundar springer genom vattnet nära en strand, med land på horisonten.
Folk tar en promenad i en mångskiftande stad.
En rad människor i röda skjortor visar numrerade plakat.
En man och en kvinna springer i ett maraton.
En person cyklar längs en gata i en ödslig stadsmiljö.
En grupp om tre löpare går förbi i ett lopp.
Bänkarna är i en lång rad med de silver runda borden i linje prydligt.
En man som sitter på ett steg.
En folksamling i en daglig rutin i en asiatisk förort.
Damen tittar på ett fönster där en stor gog slickar på läpparna.
En ung pojke klädd i smutsiga kläder ligger på en vävd matta i grunt smutsigt vatten fyllt med sopor.
Ett barn rider bak i en träkärra.
Smickrande kvinna i ett blått förkläde som står framför en hög med väskor och lådor.
En man använder en droppare för att utföra ett experiment.
Två unga pojkar, den ena håller i en påse, den andra en Unicef hink.
Två unga pojkar hämtar vatten med en unicef pail.
Två vithyade och en mörkhyad man sitter sida vid sida i jeans och svarta skjortor.
Två kvinnor står nära en grupp cyklar.
En medelålders man med mörkt hår som lagar mat och bär ett rött förkläde.
En liten flicka i röd jacka kramar en liten pojke.
En skjortlös man i blå jeans springer nerför en docka mot kameran.
En kvinna som går på trottoaren, i stan.
En man i vit skjorta och blå jeans pratar i telefon nära gatan.
En baby inlindad i filtar är instoppad i en metallvagn.
En bild av en byggnad och trottoar, människor är synliga i fjärran
Det här är torsdag kväll på lokalklubben, vänta till fredag kväll.
En man sitter i en klassisk bil medan han ler och håller i en plastmugg.
En man på gatan, stående över några konstverk, medan flera människor passerar förbi.
Två unga, blonda bröder har sina armar utspridda, den ena bakom den andra mitt i ett gräsfält.
En arbetare klädd i en ren kostym polerar en stor spegel.
En person med en blå skjorta och byxor sitter på en bänk utanför.
En tonårstjej i en rosa tanktopp med två tummar upp.
Två magdansare dansar bredvid en tegelvägg.
Kvinnor som korsar gatan framför en svart bil.
Två personer joggar tillsammans nära vattnet.
En kvinna äter en idiot utanför en byggnad.
Ett barn i röd skjorta springer runt i vatten.
En hund hoppar över ett hinder.
En prickig hund som leker på ett basebollplan med en annan hund.
Sex personer på ett möte i American Business Club.
En man i vit skjorta och röd slips pratar med folk på en restaurang.
En man i blå skjorta använder en spatel för att röra om i maten på en grill.
En man och kvinna är avbildade bakifrån sitter tätt tillsammans på en soffa medan de spelar Nintendo DS
En man spelar schack med en ung pojke.
Människor från spädbarn till äldre verkar exalterade som en kvinna i en gul skjorta hoppar ner från marken framför en skylt som säger "Bienvenue WELKOME".
Folk går runt på en karneval där stora uppstoppade djur visas upp.
Två försäljare med röda och vita paraplyer är ute i mitten av en massa människor.
Många människor i gathörnet med bruna byggnader.
Två kvinnor, en med en plack, en med namnbricka, på ett matställe.
En grupp människor i olika åldrar på en konferens pratar.
Fyra kvinnor tittar på ett fotoalbum.
En äldre man öppnar en present.
Två unga pojkar med röda flytvästar sitter bredvid varandra på däcket på en båt.
En man och en dam som båda bär vita skjortor tittar ut i fjärran.
En man som bär alla vita och solglasögon kramar en kvinna bakifrån.
En man är på en cykel framför Eddies sweetshop.
Fyra flickor spelar fotboll medan en vuxen tittar över dem.
En man och en flicka sitter på en bänk medan de äter glasstrutar.
En man i orange skjorta och baddräkt rullar i en plastboll genom vatten.
En man som fiskar under ett paraply.
Ett afrikanskt barn med en träpall på huvudet och ett annat afrikanskt barn bakom sig
Flera kvinnor sitter med ledstänger på en lutande skyttel.
En ung man som sitter i mörkret och bär en vit skjorta med handen vänd upp ansiktet med hörlurar.
En man och kvinna som tittar på grönsaker.
Tre små barn som har kul med vatten från en brandpost på trottoaren.
En asiatisk kvinna tävlar i vinterolympiaden.
En flicka klättrar på en stenvägg.
Person som går ner för upplyst tunnel med grönt ledstång.
Människor som går på en livlig gata i ett främmande land möjligen.
Två flickor sitter i lägerstolar runt en lägereld.
En medelålders man i vitt hat, marintröja och khakibyxor sätter en golfboll.
Två personer i randiga skjortor sitter vid ett bord.
Fotgängare ger efter för en brandbil när den kommer in i korsningen.
Gatumusiker spelar dragspel, fiol och gitarr.
En kvinna i vit skjorta visas bakifrån på en kyrkogård.
En man med kryckor passerar bakom en vit lastbil.
En kvinna går förbi med sitt barn och sina tillhörigheter i korgar på ryggen.
En asiatisk man som slaktar en gris som hänger på en krok.
En kinesisk konstnär och skrivare sätter upp sin skylt för visning.
En man som går med en kundvagn i en t-shirt som lyder "Långt leve de döda".
En brunhårig man med skrynkligt skägg och grön skjorta med kamera
En skateboardåkare som gör ett trick från en kvartspipa.
En man som tvättar hörnet av en jacka i en offentlig fontän.
En person går vid bron.
Massor av människor som sitter längs en låg vägg framför gräset med byggnader som kantar längs vägen.
Två män i hatt går förbi en gammal vägg.
En man i en orange turban står framför en korg med ett paket marlbororötter och andra små föremål.
En liten flicka kisar och tittar in i en lins.
På regniga gator stannar en motorcykel med två hjälmar för en vit bil.
En grupp människor går nerför en stad gata.
En kvinna i blå klänning tar en bild av en staty.
En polis i Minneapolis står framför en underklädesreklam.
Ung man i grön skjorta spela xylophone för publik i offentliga området.
En ung dam sitter i en blommig miljö med en sportdryck i handen.
En trupp i senapfärgad uniform marscherar bakom en truppledare som håller i ett svärd.
En upptagen utomhuskiosk för att sälja föremål.
En man i grönt med skägg och vit hatt går bredvid en stor orange vägg.
En rad människor för en karneval rida.
Många människor står på stora stenar som låg över en flod.
Folk simmar i vattnet nära en lång brygga.
Ett band spelar en show på kanten av vattnet på natten med en levande dansande publik.
En kvinna vid universitetet i Nottingham som leker med ett barn.
Ett amoröst par med vatten framför sig, en gammal byggnad med utsmyckade pelare i bakgrunden.
En liten flicka i rött stannar och håller en leksak i båda händerna och ler.
En grupp människor som sitter utanför ett hus med en målning av en cowboy i en röd skjorta på sidan.
En flicka i rosa skjorta klättrar upp på en trästol.
En ung pojke står bredvid en stor hög med jord.
Barn leker på en lekplats.
En man på en mobiltelefon som går förbi fyra tecken som alla säger "Aldrig sova igen"
En man går på stranden medan han bär skorna.
Två vuxna hjälper till att dela ut tårta till barn i ett klassrum.
Två unga pojkar står på en grussluttning i dagsljus.
Ung pojke i blått och ung kvinna i turkos sticker ut sina tungor för kameran.
En väggmålning av en man och kvinnor på sidan av en byggnad.
En del barn kommer ut för att leka på en gårdsplan.
Ett barn som leker på en swing set med byggnadsarbetare i bakgrunden.
Ett barn ligger på golvet och ritar en bild av en flicka, och två andra barn tittar på.
En pojke sitter ensam på botten av en stentrappa.
En närbild av en mycket upphetsad ung pojke.
En man i blå skjorta som går längs en bergsväg med getter i vägen.
En ung man ler och pekar på något utanför kameran, medan han står framför en uppvisning.
Arbetare städar upp och bygger om på en byggarbetsplats.
Två flickor plockar gula blommor en solig dag.
Två hundar leker på gräset.
Två vita hundar tittar ut på gatan och sitter bredvid en vit cykel.
En grupp människor dansar på en restaurang.
En grupp asiatiska män och en asiatisk kvinna slappnar av i en slaktarbutik.
En man som avslöjar en lastbil full av blomkrukor.
En man som sitter i närheten av högar av att producera skalning av en grönsak.
En kvinna skriver ner något medan hon väntar på ett masstransportstopp.
En man i grön skjorta och grå byxor som går på en gata och passerar förbi en affär.
En kvinna i röd klänning går nerför gatan.
Grupp av människor som har en stor kul på gatorna i sin stad med ballonger och flaggor.
Arbetstagare i gröna skjortor väntar på flera kunder.
En ung man rider en häst genom en grupp människor medan han pratar på sin mobiltelefon.
En man i rullstol sitter framför en väggmålning av en rädd kvinna.
En kvinna i ett grönt förkläde ristar kött från ett djurkadaver.
En kvinna sitter med sina blomkorgar.
En man som sitter på en pall framför ett bås som säljer fotbollssjalar.
En man med cigarett i nunnakläder.
En nunna har en cigarett i munnen.
Ett litet barn i en vagn en solig dag.
Vi ska ta det här fotot tillsammans och sätta det i ansiktsbok.
Folk pratar på en loppmarknad.
En äldre man med randig skjorta väntar på att någon ska köpa hans blommor.
Två skjortlösa män som går på en fullsatt strand.
Folk går runt på en livlig trottoar på natten.
En stor grupp cyklister rider runt på en stor bro.
Dussintals cyklister cyklar på en hängbro utan synliga bilar.
Det finns en grupp unga män som är hopsnärjda i en cirkel, till synes sjungande.
En man i en blå jacka med vita byxor står utanför en röd tegelbyggnad nära en annan man som håller två gula väskor.
Folk passerar signalen.
En liten asiatisk pojke går nerför gatan i traditionella asiatiska kläder tittar tillbaka på en dam klädd i höga klackar och en beige kjol.
En man står framför en grönsaksutställning.
Asiatisk gatuscen med två kvinnor i förgrunden, röd byggnad med lejonaffisch i bakgrunden.
Fyra tonåringar hoppar med bollar på en basketplan.
En man med lila skjorta, blå gympaskor och en svart ryggsäck som cyklar.
En mörkhårig kvinna som går medan hon håller sitt barn.
En brun hund som bär krage jagar och biter på en röd kvast.
En grön bil parkerad nära ett trångt utrymme.
Två män i en by i Indien spelar pinneboll.
Vissa människor går på gatan nära en mycket stor väggmålning.
En grupp musiker som spelar musik framför en byggnad.
En man som håller färska frukter framför en marknad.
Grupper av turister går över bron och tittar på utsikten över gamla byggnader.
En leende kvinna med svart smet över ansiktet håller i ett paraply.
En clown i vit skjorta och slips som spelar fiol.
Två kvinnor i en grupp ler tillsammans.
En man som bär bast och tonade glasögon står framför en mikrofon.
Fotgängare går på trottoaren i en urban miljö.
Ung flicka med kort, mörkt hår bär en rosa skjorta klättra trappor framför cyklar.
Tjejen sticker ut tungan medan hon hula hänger med två korgar
En svart manlig idrottsman som gör ett hopp under en tävling.
Ett par campar i skogen.
En kvinna i blått bär glasögon håller upp en blå och vit randig skjorta till en pojke klädd i gult som också har glasögon.
En hund bär ett gult rep över klippor som är täckta av sjögräs.
En man i kostym sitter utomhus och använder sin bärbara dator.
Fem personer står på gräs.
En kvinna med röda skor står mitt på gatan.
En man som fiskar i vatten med stora vågor.
En kvinna som pratar i telefon bakom ett rack med de stora blå plastflaskorna.
En man tar ett foto i fotots riktning.
En man sitter nära en annan man som står på trottoaren.
En publik sitter på en veranda utanför.
En man på scenen visar sitt kökort för sin vän.
En man med röd skjorta och svart hatt stirrar på en annan man.
De tre männen leker med en frisbee.
En pojke och flicka kysser varandra vid en sjö.
En man som sitter på en stol med benen korsade och tittar åt höger.
En man på en hiss inspekterar fasaden på en byggnad.
En man och en svart väst som dansar med en kvinna med svart hår.
En fågel-ögonblicksbild av människor som står runt och håller sina drinkar.
En kvinna och en man och ett barn står på en gata med paraplyer
Två personer bär röda hoodies rider sina cyklar nerför gatan.
Ett par omfamnar mot en grövre pelare medan en man fotograferar.
Två män handlar på en upptagen asiatisk marknadsplats.
En man i blå skjorta går mellan klippor i grunt vatten nära en naturskön tropisk strand.
En ung man som bär jeans balanserar på ett tågspår.
En person som sätter upp sitt hår i ett livligt område i en stad med flera telefonkiosker i bakgrunden.
En man som sitter vid ett vitt plastbord i skuggorna.
Killar och flickor på ett trångt ställe med drinkar i handen.
Två barn står med ett nät vid en grunt strand.
En kvinna med solglasögon jobbar med en kontrollbräda.
Flera människor står runt på en fest.
En grupp människor pratar med varandra i en bar.
En man sitter i en stol på gatan och spelar gitarr.
Två män med fiskespön står på en strand
En fotbollsspelare i grönt tar itu med en fotbollsspelare i vitt.
En man i blå jacka och vit hatt poserar med en gammaldags kamera.
En man cyklar förbi en orange vägg utanför.
En grupp människor som rider på ett promenadbälte på flygplatsen.
Folk står på trottoaren på en gata.
En kvinna får mat under ett blått tält.
En grupp unga dansare uppträder tillsammans framför Radio City.
En grupp dansare uppträder med matchande kläder.
En man skateboardar förbi en graffititäckt vägg.
En kvinna står och tittar ut över vattnet medan någon tar en bild
2 våta pojkar i blå baddräkter
En gammal man sover i en stol utanför en övergiven byggnad.
En svart kvinna som sitter med en asiatisk flicka med falska tatueringar.
En man sitter i en stol och spelar gitarr.
En kvinna som tweaking något på en cykel hängande från ett staket.
En man med röd hatt, röd jacka och röda solglasögon lyssnar på sin musikspelare.
Tomten är i linje med dansarna för paraden.
En kille som bär en blå jersey #5 träffar en gul softball i ett gräsfält till några fältare.
En brun katt sitter ovanpå en gammal bil.
Man och kvinnor sitter på trappan på kvällen med många pelare runt dem.
En vit katt sitter på en vägg.
En man som bär svart jacka och hatt går och håller i en cigarett.
En kvinna med sitt barn väntar på en bänk.
En ung kvinna sitter på en röd buss och tittar ut genom fönstret.
Dussintals människor går på ett stort torg framför en massiv trappa.
En ung man som tar bilder när andra civila går förbi honom.
En man använder en kamera på en stadion.
En man i svart jacka står bredvid en väg som har utsikt över en vattenförekomst.
Folk klädda i gröna uniformer plockar upp metall.
Två män sitter vid ett bord med drinkar och tittar på en annan man som går med en väska.
Folk går och en kvinna bär väskor.
En kvinna med blå skjorta, jeans och röda konverserade gympaskor tar ett fotografi.
Utsikt över den historiska delen av en europeisk stad.
En kvinna klädd i blått och bär solhatt ler.
En asiatisk kvinna som står i ett trångt stadsområde och lyssnar på musik.
En man som cyklar försöker korsa en livlig gata.
Ung pojke i svart skjorta sitter på mödrar axlar
En kvinna (Carol Thorn) i en röd klänning som spelar en elektrisk cello på en scen.
Folk som sitter på en uppsättning blekmedel.
Tre män sitter på ett steg bredvid varandra.
En utomhusförsäljare med ett bord fullt av hattar, dockor och smycken.
Två munkar i orange rock talar utanför ett hus där en man i normala kläder går ut.
Kvinnan leker med ett barn.
En man i vit skjorta och khakibyxor passerar framför ett mellanmål.
En grupp äldre män sitter på en bänk inomhus.
En kvinna som bär en röd klänning spelar ett stränginstrument.
En del människor står i en stor grupp av hjul.
Flera människor samlas vid ett parasoll toppade bord strax utanför en butik som heter DAHLAK.
En person har två små barn som sitter framför honom på en motorcykel.
En man håller upp den vita skjortan han bär exponerande är buken medan han sitter på en röd motorcykel.
En asiatisk kvinna håller sitt barn, som bär en blommig jacka.
En militär marschtrupp av soldater i formell uniform med röda rockar och luddiga svarta hattar marscherar förbi, ledd av saxofonisten.
En man ryser med sin kamera.
En kvinna med kort hår spelar fiol.
En flintskallig man med glasögon och en svart skjorta som hullar ett instrument.
Ett par står högst upp på en trappa utomhus och kysser varandra.
Mannen i den blå skjortan cyklar nerför gatan.
En man klädd i kockkläder som håller en stor sked över en stor gryta på spisen.
En mycket upptagen gata sida med många människor interagerar tillsammans nära en kinesisk restaurang.
Flera motorcyklister rider längs vägen en solig dag.
Ett par turister på en kinesisk marknad tittar på sin kamera.
En ung modell poserar för sin fotografering under en docka.
En flicka går förbi ett fönster med en handväska.
En familj står på en tegelgata och pratar med en konstnär som håller i en stor skissdyna.
Folk går genom en gränd i Turkiet.
En liten skara människor samlades för att titta på verksamhet som inträffade framför dem.
En kvinna i blå jacka går längs en väg.
En person klädd i svart med en röd ryggsäck som går mot en utomhusmarknad.
En färgstarkrickshaw med två beskyddare på stranden som stannar vid en kokskiosk.
Tre män kikar genom ett stängsel som är täckt av stenar.
En man verkar spela något slags instrument.
En pojke som bär röda badbyxor svingar från ett rep ner i vattnet.
Gatuförsäljare i Europa säljer till flera äldre.
Tre män klädda i blå spela gitarr medan en kvinna sjunger.
Ett band spelar en spelning för en publik.
Ett band spelar på scen med två personer som står vända mot varandra och sjunger, en person som spelar trummor, en på tangentbordet och en person på gitarr.
Ett jazzomslagsband spelar under heta strobeljus.
En person går nerför en korridor av sten valvbanor.
En brud på sin bröllopsdag bär sitt orange bälte.
Kvinnor i en vit skjorta med en halsduk som går medan hon sms:ar på sin telefon.
En blondhårig kvinna i en benvit kappa skjuter fåglar från ett bord.
En afrikansk amerikansk pojke står i en bur med handen mot ansiktet.
En flicka står i närheten medan en pojke sitter i en öppen dörr.
En grupp människor slutför ett drag med huvudet något sänkt och armarna böjda och upp.
Tre personer går framför en mycket reflekterande byggnad.
Två kvinnor bär solglasögon och äter mat.
En skara människor samlas i ett gräsbevuxen område.
Kvinnliga vakter står i en grupp med solglasögon på.
Man i svart skjorta rider kollektivtrafik.
En vy nerför en stadsgata från ett parkcentrum.
Skotska män i formell klädsel spelar säckpipan.
Folk är uppradade mot varandra med flaskor med bärnstensvätska, lådor och etiketter.
En mörkhyad man framför en vibrerande röd, svart och vit bakgrund.
Två personer kysser varandra på en mycket utsmyckad balkong bredvid stora pelare.
En äldre man med käpp är ute och handlar.
En man i vit skjorta tar betalt för mat från två kvinnor.
Fyra äldre män sitter ute i stolar.
En stor grupp människor går utanför förbi en McDonalds.
Flera människor går ut i regnet.
En man står framför en vit vägg med en företagsannons på sig.
En skara människor som sitter på en gräsmatta klappar.
Det finns rosa konstgjorda tulpaner i ett matställe, med tre personer i bakgrunden.
En arbetare i spritbutiken.
En man i grön skjorta klipper gräset i en gräsklippare.
Fyra personer avbildas i en katedralliknande byggnad.
En kvinna med kort brunt hår, i jeans och en leopardtopp tar en bild.
En man utan tröja som sitter på en moped.
En kvinna som bär en blå t-shirt som säger Nike och bär en grönsak.
En kvinna i randig skjorta visas ett halsband.
Två kvinnor i shorts sitter på trappan till en lägenhet eller hus.
Folk flyttar hemifrån.
Den orangehåriga hunden skakade på huvudet medan han stod på stranden.
Medelålders man med långt blont hår och glasögon sitter med en publik.
Ett ungt par som pratar med en äldre kvinna på en livlig plattform.
Ett barn som står framför en gigantisk mekanisk elefant.
En kvinna hjälper en flicka att rita en symbol i stenarna.
2 kvinna går nerför gatan bredvid graffiti
Två motorcyklister rider nerför en gata.
Ett par barn sitter på en bänk och leker med en röd hjälm.
En man sitter utanför sin korvkiosk bredvid en byggarbetsplats medan han läser en bok.
En grupp människor låg i parken.
En man och en kvinna stannar för att ta en bild i en utomhusmiljö.
En man i en blå jacka pratar in i en mikrofon.
En man i svart t-shirt och svarta shorts dammsuger i ett sovrum.
En flicka i parken tar en bild.
En liten pojke som krattar löven med en kratta.
En liten asiatisk flicka står på gatan och håller i en röd väska.
Paren dansar på gatorna.
En man står bredvid en stor svart lejonstaty.
En kvinna i svarta byxor korsar en livlig trottoar framför en herrklubb.
Åskådare tar bilder på en cykeltävling.
Mannen leder sin svarta och vita hund över ett blått hinder.
En man beställer en korv från en gatuförsäljare.
En ung blond flicka håller en strandboll mitt på ett gräsfält.
Tre unga flickor går nerför en trottoar.
En grupp pojkar går genom en plaza.
En man sitter på en kedja.
En kvinna som står mot en byggnad och tittar på sin telefon, med benet uppstött.
En ung man kollar sin telefon medan han lutar sig mot en tidningskorg.
En ung man utan tröja står nära en bil med surfingbrädor på sig.
En kvinna som bär en avtrycksrock läser en bok.
En man går nerför en gata där husen är målade i ett geometriskt mönster.
Bilar och motorcyklister kör nerför en gata kantad av gamla byggnader.
En stad gata med frukt vagnar och en buss, och massor av människor.
En man i vitt sitter utanför med en kattvän.
En kvinna i blå topp och solbränna målar ett barn kramande träd.
Två arbetare arbetar med ett verktyg och fäster ett föremål i sten.
Folk står på gatan utanför några höga gräddfärgade byggnader.
En busker uppträder på gitarr bland en fullsatt gata.
Sju flickor står i kö för att spela i parken
Två kvinnor klädda i vitt står på trottoaren under ett paraply.
Man i khaki byxor böjd över framför en vägg täckt av graffiti.
En skjortlös blond man spray målar graffiti på en vägg.
En kvinna i vit skjorta och Jean shorts står med en dryck i vänster hand.
En man på gatan spelar trummor på gamla burkar.
En kvinna i allt rosa och guld stirrar på något.
Folk samlades utanför en kyrka i trappan.
En man med en portfölj som gick i ett område målades på väggar.
En ung man lyssnar på hörlurar på gatan.
En kvinna som står på en korsning som bara har handen och långfingret lyst upp.
En kvinna står i en pool med tre unga pojkar.
En dam simmar med två unga pojkar som båda bär gröna vattenvingar.
Två män i hattar som gräver upp stenar och jord.
Tre flickor med långt brunt hår sitter bredvid varandra nära ett träd.
En ung kvinna går genom sittande åskådare.
En kvinna med svart pennkjol och vit knapp-up skjorta med flip-flops går tvärs över gatan.
Två personer sitter på sidan av vägen framför en karneval.
Två asiatiska män med hårda hattar på en röd skoter passerar av två människor som knäböjer på vägen med två korgar på sidorna.
En pojke ger "tummarna upp" medan vattenskidor på grumligt vatten.
En ung man fotograferar två vänner bredvid havet.
En man med långt skägg tittar på vattnet.
En man breakdancing på en stor matta medan vissa människor tittar.
En grupp ungdomar som väntar på att gå över en gata.
En man i svart skjorta och vita shorts breakdances framför åskådare.
En cyklist rider ensam i ett avlägset område hoppa över objekt.
En ung flicka i glasögon observerar något i fjärran.
En person i rosa vattenglasögon blåser bubblor under vattnet.
En kvinna i klänning i solglasögon och en man i blå skjorta står utanför med en stor publik.
En kvinna bär blå shorts, en gul blus och solglasögon.
Två flickor står vid vägkanten.
Denna cykel hoppa verkar sätta skyline i anslutning till ryttaren.
En man i vit skjorta vandrar över klippor och vatten.
Tre bruna valpar springer i gräset.
Två personer plockar upp sina tillhörigheter framför en Subway.
En skäggig man fotograferar med kamera och lång lins.
En man som bär glasögon sitter framför en Apple-dator och dricker ur en kopp medan en annan man som bär mössa och glasögon står framför en mikrofon.
Män sitter på påsar på marken.
En man klipper håret på en öppen plats.
Tre killar som hänger utanför ett fruktstånd.
En baby som hänger i en hoppare på ett däck vid en hamn.
Barnen går nerför gatan bredvid biltrafiken.
Tre män badar i en kanal utan sina skjortor.
Några barn som spelar tv-spel.
En dam i röd skjorta och bikini nedredelar är på väg att surfa på en blå bräda i havet.
En soldat pratar inför flera människor.
Folk är på en berg-och dalbana framför en vattenförekomst.
Man och kvinna tittar på en lott i Kina.
En ung, skjortlös pojke framför en pool medan en kvinna i religiös klädsel står bakom honom.
Damen spelar en omgång hopscotch.
En kvinna med gul hatt och flerfärgad klänning undersöker en bok på en uteplats.
En person och ett barn rider en gräsklippare nerför vägen.
Mannen i gul skjorta tittar in i sin blå tvättväska, bredvid en tvättmaskin.
En man som driver tunga maskiner.
Mannen i den grå skjortan blockerar den andra personen i den svarta skjortan ur sikte medan han tittar in i tvättmaskinen.
Två äldre kvinnor går i grunt vatten.
En äldre blond kvinna med solglasögon som lutar sig mot ett broräcke en solig dag.
En hemlös man sitter och stirrar
Heavyset kvinnor i en blå och vit klänning går nerför ett kvarter.
Tre vänner som hänger i ett fotobås.
Två män skrattar framför ett ljus.
En flicka sitter mot en byggnad nära en brandpost.
En svart man sitter vid ett bord och fotograferar en äldre kvinna på en uteplats.
Två kvinnliga poledanser mitt på gatan.
En man försöker ta en bild av en kvinna och sig själv kyssas medan de står omgiven av blommor.
En gentleman som sitter ensam vid ett bord.
En person som bar gråa konverserade skor tog en bild av vattnet och rörde knappt vid skorna.
En grupp män klädda i konstiga kläder talar om sin dag.
En kvinna och man vid ett skrivbord med massor av kontanter eller valuta runt dem.
Gnistor flyger som en man svetsar stål.
2 män och en kvinna som bär rött håller en surfbräda stående i sanden.
En del barn leker i gräset utanför nära ett träd.
Två kvinnor tittar på åsnor på en strand.
En grupp människor står längs stranden.
Två män leker med sina svarta och vita hundar på stranden.
Två gamla män sitter på en parkbänk.
En kvinna med grön handväska sitter på en bar med ett tomt glas framför sig.
En bartender förbereder många blandade drycker.
Kvinnan i en svart baddräkt, som ligger på en säng, ovanpå en byggnad, med ett högt vitt paraply inom synhåll.
Två kvinnor skrattar åt ett skämt på en stoppskylt.
En pojke i röd skjorta med ett rött hjärta rakat i sitt blekta hår pratar på en mobiltelefon.
En man med röd skjorta och jeans som går genom ett centrum.
En asiatisk fotograf kollar sin kamera framför en modebutik med fotgängare som går runt honom.
En person som surfar på vågens krön.
En man med stort vitt skägg knuffar en vagn full av sopsäckar och kartong nerför en trottoar.
En man som spelar trummor på upp och ner kannor.
En gammal person tittar på TV medan han sitter på huk framför en butiksdisplay.
En man i en blå t-shirt och en ansiktsmask arbetar med krokar.
Två personer simmar i en stor pool som omger av strandstolar.
Två reparatörer i hårda hattar arbetar på en byggarbetsplats.
De flesta av dem bär mask för att skydda dem från föroreningar.
En flicka springer på gräset.
Två barn rider på baksidan av en trehjulig scooter som drivs av en ung dam i rosa.
En byggnad har ett bi målat på taket.
Blonda barn sover på ett vuxna knä när de åker buss.
En kvinna i klänning, som håller ett uppstoppat djur, handväska och paraply, stående i regnet.
En kvinna ger kameran ett smutsigt utseende när hon går nerför trottoaren.
Två personer med stora öronproppar sitter bredvid varandra.
En svart kvinna med en halsduk på huvudet står på en trottoar och ler.
En ung dam går på gatan.
Två män rider på en motorcykel på en väg.
En kvinna äter popcorn från sitt popcornstånd.
En kvinna ute på gatorna i en svart skjorta som pratar i telefon.
Ett stort antal äldre människor sitter på bänkar utomhus.
Folk i affärskläder, gå längs en gränd.
En sfärisk formad havsakvarium byggnad.
En man sitter i en Exuma med tre andra män som står runt en byggarbetsplats.
En blond kvinna som bär en tank topp och olika färgade handskar.
Flera ungdomar spelar ett brädspel med hjälp av en stor filt i ett gräsfält.
Två personer går och tittar på uppstoppade djur.
En grupp människor tittar på böcker i ett bibliotek.
En kvinna läser med ett barn.
Ett gäng kvinnor i ett bibliotek med barn.
Människor som går på en asfalterad gångväg nära en hamn.
En äldre gentleman sitter på en bänk och röker en cigarr med korsade ben.
En livlig utomhuspark i Europa.
En kvinna i blå kjol som knuffar en barnvagn längs en trädkantad gata.
En volleybollspelare som slår till mot en volleyboll.
Mannen i vit skjorta och mörka byxor lutar sig mot en vägg med två skyltfönster som har starkt ljus.
En man i grön hatt och randig skjorta som går.
En kvinnlig motorcyklist med hjälm i handen står vid sin cykel.
En kvinna med grön väska tar en bild.
En kille i svart skjorta och bruna byxor lutar sig lite ut genom ett stort fönster och tittar på något.
Ett ungt par som kysser vid en cykelrake.
En man som målar framför en butiksvägg, hans målningar visas.
En man pratar på sin mobil framför en fontän.
En flicka är i luften framför någon form av kalistik eller kanske dyka ner i en pool.
En gymnast i svart och orange kostym i luften.
En dam med svart hår och en vinröd och svart kostym utför ett dyk.
En man som tvättar fönster på en röd tegelbyggnad.
En ung kvinna som bär en glittrig svart kostym glider över isen.
Folk tittar upp på ett flygplan som flyger förbi
En man i vit skjorta talar med en grupp på sju barn.
En äldre man med vilt hår kollar in motorcyklar.
En kvinna i röd rock sitter i gräset med kaniner.
Ungefär sex äldre kvinnor sitter på en bänk och pratar.
En afrikansk man i en färgglad hatt spelar kongotrummor.
En man som bär en gul hatt drar i ett rep.
En grupp män i smoking pratar med folk som sitter på trottoaren.
En ung kvinnlig simmare får en tröstande kram från en tränare.
Ett vackert gatufoto där människor går förbi en gammal byggnad.
En kvinna och gamla damer sitter på en bänk
En pappa och en son njuter av en cykeltur på en solig dag.
Attraktiv kvinna i svart med sin mobiltelefon.
En kille i svart baddräkt som kliver ur poolen på ett hotell.
Man står på fotboll med knän medan två kvinnor tittar.
En liten flicka med en gul skjorta som hoppar över en orange kon.
En ung flicka som hoppar över apelsinkottar.
En äldre man i en orange ceremoniell jacka har en massa blommor.
En man i blå skjorta bär en väska över sin högra axel.
En ung person med dekorativ ansiktsfärg som liknar en tigers markeringar snarrar.
Flera löpare tävlar i en road race.
En liten flicka gör ett handstånd medan hon ler
Kvinnor som cyklar på en gata.
En kvinna med en vit handväska går över en grå plattform framför en hög byggnad.
En man bär clownmakeup.
En man med bruna byxor säljer mat från en mobil automatgrill.
En man har lite pappersarbete om bankräddning.
Ett barn som bär en röd skjorta rullar en bowlingboll nerför en fil.
En kvinna med en designväska beundrar utsikten.
En man cyklar förbi Chung May Food Market.
En affär är öppen på natten.
En man i tung makeup och en blodig skjorta håller i en vattenflaska.
Folk cyklar i en allmän gångväg.
Cyklare deltar i en tvåvägs street ride, med banor åtskilda av gula kottar.
Två bilar tvättas på en parkeringsplats.
En pojke med jeansshorts och ljusblå sneakers rider en skateboard bredvid ett högt staket.
En ung kvinna klädd i svart tittar på artiklar från en gatuförsäljare.
En tonårspojke med röd hatt sitter vid sidan av en gångbro medan människor går förbi.
Folk i ett matställe som skrattar och pratar.
En solig dag är den här tatuerade mannen klädd i en detaljaffär.
En livlig stad med bilar och människor med en jättestor skyskrapa.
En grupp amerikanska kamelryttare på en grusväg som ler och har kul.
En blond kvinna som håller något i handen medan en annan kvinna och man går förbi henne.
En man som läser en bok på trottoaren med bara sin blå pyjamas och hörlurar medan han sitter på en stol.
En cyklist med barn i ett litet fack med cyklister i bakgrunden.
Ett barn i en jeansjacka med "Kärlek dödar långsamt" skrivet på baksidan av den.
Folk går på gatan medan andra sitter och äter lunch.
En fotbollsspelare lägger ner skadade som assisteras av domaren och en annan spelare.
Två män bär nät nära en pier.
Två kvinnor leker i vattnet på en strand nära strandlinjen.
En grön halvtäckt bro finns framför ett hus.
En liten flicka i en gul t-shirt tumlar mot slutet av en gul rutschkana.
Tre personer, alla klädda i mörka kläder, står och pratar i ett gathörn.
Dinosaurieutställningen ligger bredvid ett träd som har en ballong fast i sina grenar.
En kille i blå skjorta drar något.
En byggnad med en stor skylt som lyder: "Smärta är tillfällig, Att sluta varar för evigt".
En stor skara står framför en upptagen byggnad.
Ett barn i grön jacka och blå hatt sitter på en bänk och äter glass ur en kopp.
Det här är en professionell dykare.
En kvinna i röd och blå skjorta stirrar på en affisch på väggen.
Två män roar sig i en skatepark, den ena cyklar medan den andra åker skateboard.
En kvinna i en grön skjorta talar på en mobiltelefon medan hon går förbi en man i en blå skjorta som sitter och läser en tidning.
Tre personer klädde upp sig och spelade musik på en trottoar.
Tre yngre män dansar framför en halvomringad publik.
Ett par elever låg bredvid varandra i en betongpark.
En man i grått och svart spelar en svart akustisk gitarr med en något kortare kvinna som bär rosa och spelar violin.
En man som utför breakdancing utanför inför en folkmassa.
En kvinna med tatueringar som bär en svart tanktopp tittar på marken.
Man i ett fält tar ett fotografi som ser nedförsbacke.
En kvinna som kör en blå cykel bär en vit stol på halsen.
En man kittlar ett litet barn framför ett soligt fönster.
En geisha står utanför en butik och kikar till sin sida.
Folk rider på en motorcykel på en strandgata.
Mannen i långärmad t-shirt sitter vid ett köksbord och äter från en pappersplatta.
En asiatisk man i glasögon och en blå klänningskjorta ger en presentation med hjälp av en projektor.
En man och en kvinna går förbi en butik.
En man och kvinna lägger handdukar på stranden.
Gatulampan är brännpunkten, men det finns en person som böjs ner direkt bakom lampan.
En liten flicka springer nerför en stig i en japansk trädgård.
En man med ryggsäck läser en bok nära en kvinna som slappnar av på en betongplatta.
En äldre gentlemän städar baren medan en man bakom observerar.
En kvinnlig artist på en scen med mikrofon.
En tågstation plattform klockan 11:27 på morgonen.
En man med blommor som tittar ut genom sitt andra storyfönster.
Kvinnan sitter ovanpå en rad block.
En schizofren man målar en karikatyr av två män trots att det bara finns en kvinna.
En kvinna fokuserar sin digitala kamera på stora evenemang.
En kvinna har ett svart paraply och en vit shoppingväska i regnet.
Människor med paraplyer går förbi affärer i regnet.
Ett par stannar på en brud för att titta på en damm.
En äldre man utför reparationer på en ung mans cykel.
En kvinna och en man sitter på en stenbänk, med höga byggnader bakom sig.
En person kryper under en filt medan han sitter på en bänk.
Två gräsklippare skär ner palmträdsgrenar i ett närliggande community college under en blåsig dag
Folk som sitter i en upptagen metropol.
En man i en flygplats vågor vid kameran.
Regn utanför och tre svarta paraplyer och ett gult och rosa paraply.
En kvinna sitter bredvid ett blomsterstånd framför en McDonald's restaurang.
En individ som trycker ner regnet från taktopparna.
En grupp människor på ett blomsterstånd ser ut som en stor mängd vattenfall ovanför tältet.
Två personer bär ryggsäckar går längs sidan en byggnad.
En person i en grön och vit skjorta rider en smutscykel nära en grupp träd.
En liten pojke springer genom gräset med en flagga.
Ett svart barn som sitter på en leksak som biter i fingrarna.
En kvinna på sjukhuset håller sitt barn
En man i blå hjälm går bredvid rök och en röd lastbil.
En gul burk i New York.
En man i stamdräkt går nerför gatan medan åskådare står bakom röd och vit barriärbyråkrati.
En kvinna i orange skjorta njuter av mat i en offentlig miljö.
Hunden med alla bekvämligheter i hemmet och ändå har inget hem.
Folk som åker rulltrappa hellre än tar trapporna.
Flera glas och keramiska föremål arrangeras på hyllor med spegelbaksida.
En kvinna läser sin bok i en lokal stadspark.
En kvinna i brunt håller sitt barn framför en asiatisk-inspirerad byggnad.
Människor som tittar på dyr utrustning och ler
En man i svart keps sitter på en bänk.
Mannen bär orange framför damm och skräp.
En skateboardare utför ett flygtrick bland dingiga väggar med kraftledningar som korsar bakgrunden.
Några asiatiska tonåringar tar ut pengar från en bankomat.
Två män och en kvinna i kostym går nerför en gata.
Två män och en kvinna står framför en spis.
En man såg mycket liten ut, när han gick längs den gamla byggnaden.
Olika människor som hänger utanför en byggnad.
En man i en grädde blazer och fedora spelar saxofon.
En person i röd skjorta och svarta byxor böjde sig över.
En kvinna i militäruniform med håret bakbundet.
Byggarbete på en väg i centrum.
Två kvinnor som bär stövlar och håller i väskor pratar med varandra.
En indisk kvinna i traditionell dräkt går förbi med ett paraply.
Denna stig leder upp till äppelmarknadens ingång.
En man som sitter på några trappsteg på en trottoar av affärer.
En man med ryggsäck som stirrar på kameran på en gul abstrakt bakgrund
Folk som kör en gammal kärra.
Två kvinnor läser en affisch på Berlinmuren
En svart bil passerar en Walgreens.
Tre män bestämmer sig för att äta en kyckling från en lokal butik.
Tre kvinnor klädda i vitt går tillsammans.
En kvinna på en scooter med en cigarett hängande ur munnen.
Den lilla flickan leker längs strandlinjen när måsen passerar förbi.
En kvinna i rött som sitter och väntar på att få sin förmögenhet berättad på en spåman.
En person i gul skjorta cyklar förbi en historisk byggnad.
Två män rakar sig vid en diskbänk när en kvinna ser på.
Unga svarta män som spelar basket i en gymmiljö.
En man går nerför en trottoar och trycker på en låda.
En upptagen, rekreationsstig nära en vattenväg rymmer vandrare och cyklister.
En liten pojke i brun och orange skjorta sitter vid en gata.
En man och kvinna tittar på många bollar på marken.
En kvinna går på en trottoar tvärs över gatan från en Discount mat- och klädaffär.
Två kvinnor drar resväskor längs en bred trottoar.
Män som kastar tomater från en stor soptunna.
Kvinnan pratar i sin telefon när hon plockar upp burritos.
Någon bär svart skjorta och shorts och en annan bär grå topp och jeans kjolar går sina hundar.
En grön Animaniac-mugg bredvid en man som skriver på ett skrivbord.
En ung kvinna som bär en svart och röd randig skjorta står framför en mikrofon, tvärs över scenen från en gitarrist.
En man och kvinna sitter på en bänk vänd mot en affisch av en kvinna.
Ett barn som saknar en sko sitter på en röd kudde.
Den här unge asiatiske mannen vilar en kort stund utanför en kontorsbyggnad.
En man som bär blå skjorta är på trottoaren och ger en annan man en skoputsning.
Folk kastar tomater på varandra.
En kvinna har en grön och vit jacka upplyft över huvudet.
En flicka knäböjer framför kanten av en klippa
En naken man som sitter i parken nära sin cykel och läser tidningen.
En kvinna täcker sitt huvud medan hon är ute i det klara solljuset.
Två små killar sitter på en tegelvägg, den yngre läser något för den äldre.
Identiska fabriksarbetare är uppmärksamma.
En blond tjej i rosa tröja håller i ett barn.
En man i bruna skor sitter mot en grå vägg.
Två stora hundar leker tillsammans på en gård med ett högt staket.
En man blåser vatten ur en pipa.
Ett utomhusevenemang med en kille som säkrar en presenning till ett skyddsrum.
En parad av något slag äger rum.
En skara män klädda som japanska samurajer slår på olika poser.
Folk går nerför en gata under en regnig dag.
En man klädd i en vit superhjältedräkt med en guldstjärna hoppar upp i luften på ett torg.
En glasblåsare gör ett vackert konstverk i sin eld.
En ung pojke med röd skjorta och jeans står mitt i ett fält och kastar ett leksaksplan i luften.
Grönt tygmaterial framför en gata, med människor som går förbi i bakgrunden.
En man i grön skjorta bär en korg över huvudet medan han talar med en grupp människor.
En cykelbud som går i parken.
En man kollar sin mobil, medan två andra män köper öl i en affär.
Olympianernas parad trängs på stadion.
En svart man utan skjorta håller i två kaukasiska blondiner, medan en flicka håller huvudet i hennes händer.
Paddlare hamnar i en vattenstrid.
En fin väg och gångväg vid en flod som leder upp till en bro.
En kvinna som går nerför gatan i regnet.
En ung flicka är ute och tittar på klänningar.
Mannen går genom ett fält och bär hö.
En grupp människor i clownmakeup uppträder på gatan.
En handikappad kvinna som spelar sport.
En asiatisk man står på en trottoar framför en röd skoter.
Två personer i smink ger ut papper på gatan.
En grupp människor med målade ansikten står utanför.
Två kvinnor som läser medan de sitter på bänken.
Två män i rutiga skjortor rider på hästar och de lassoar en kalv.
Folk spelar sport och bär gröna skjortor.
En vit man sitter på en brun häst när han svänger en lasso runt ovanför huvudet.
Två pojkar med gröna skjortor som spelar pingis i en turnering.
En äldre man, en medelålders man och en ung man sitter var och en på en häst och tittar åt olika håll, i en fålla nära ett stort träd.
De två männen rider på hästar för att jaga en vit häst.
En medelålders man i Supermanskjorta och knästrumpor går nerför en trottoar förbi en tegelbyggnad.
En ung flicka blåser fröna av en maskros.
En kvinna som rider en brun och vit häst som försöker repa en kalv.
En man i cowboyhatt rider en brun häst.
Man leder en kohjord nerför en stig medan man rider på en häst.
En cowboy bär en brun skjorta som säger att USA:s armé håller i en hästblya.
Två män rider på hästar och pratar medan andra män också rider runt dem.
En liten pojke som leker på en lekplats.
Tre kvinnor och en man sitter i ett rum med två instrument.
En man som spelar på vägen och en boll springer.
En man på hästryggen, inne i en inhägnad, jagar en stut.
Ett par väntar nära sina väskor, när några vandrare passerar.
En kvinna i en rosa tanktopp rider en häst i en rodeo.
Två ryttare jagar en ko runt på tomten.
En kvinna i bikini övredelen som har en tatuering på ryggen tittar åt vänster.
En kvinna som rider på en häst slår en ko.
En person som rider på en häst och försöker repa en kalv som springer från dem.
Två killar en kille jag befriar en vit häst.
Två kvinnor går nerför en trottoar, en bär svart skjorta med röda byxor andra bär blå tröja med jeans.
En kvinna repar en kalv i en rodeo.
En man i orange och vit randig skjorta som sitter på en båt och pratar i telefon.
En mycket lugn, fridfull sjö med ett berg i bakgrunden och en man som fiskar.
En man i gul skjorta som står vid ett långt bord och tittar på olika sorters blomsterarrangemang på bordet.
En grupp tittar på saker till salu.
Många skjortlösa och stökiga män spelar ett spel.
En mörkhårig kvinna med röd kjol och vit topp använder en telefonautomat.
Tre barn leker på gräset under ett mångfärgat paraply och bär regnbågsfärgade kläder.
Några går nerför en gata.
En brud pratar med män på sitt bröllop.
En liten hund som bär en denim minikjol.
En ung flicka som håller i ett litet barn som bär blå overall.
En man rider gömde Rickshaw på en övergiven gata.
En flicka n en orange klänning rider en cykel på en annars tom gata.
En grupp motorcyklister rider nerför gatan.
En äldre asiatisk man sitter på stentrappor i vad som ser ut att vara en affärsmiljö i centrum.
En man i svart tröja går tre små hundar.
En man i svart skjorta tittar på kameran; olika textilier kan ses hängande i bakgrunden.
En kvinna på en skoter stannar vid en stadskorsning.
En man utan skjorta på att gå bakom en maroon Ford lastbil.
En man med lei är runt halsen och håller i en mikrofon.
En man i blå skjorta går över en bro.
Bilar parkerar i en närbutik.
Många sitter vid ett bord med gröna paraplyer på.
En man utan tröja som går bakom en lastbil.
En äldre kvinna som knuffar en vagn fylld med lådor går vid teaterskylten mot "South Pacific".
En kvinna i svart skjorta med gult pannband sitter med kaffe.
Tre personer inklusive en långhårig flicka med uträckt arm och handflata upp.
En person som står utanför en gammal byggnad med hörlurar på.
En man i svart hatt håller en mobiltelefon framför ansiktet.
Ett barn leker i en Wiggles bil medan en man tittar.
En äldre man tittar på en kvinna i gul skjorta medan de sitter på bänkar framför en sten- och gipsvägg.
En man i blå skjorta pratar i telefon.
En kvinna med solglasögon går förbi en tegelbyggnad i staden och kollar sin mobil.
En kvinna i svart skjorta tittar på sin kamera.
En man i svart läderjacka som vänder ryggen till en soptunna.
Män i vita kostymer står i vägen och längs sidan av vägen.
Två personer, en i röd skjorta, sitter vid vattnet mot några båtar.
En man och kvinna står med två röda cyklar.
En äldre man med sin hårda hatt i handen, står och stirrar på något.
En man på en cykel rider genom en liten publik.
En man, med en hund, håller i koppel och en liten väska.
Det här fotot finns i ett annat land, som Japan?
En man som spelar ett instrument under några trappor och en röd bil i bakgrunden.
Paret slappnar av på trappan och studerar guideboken.
En man och ett par kvinnor förbereder ett gult fordon med förnödenheter att ta till en destination.
En kvinna pratar med en man.
En man och två kvinnor är nedlåtande en säljare på gatan.
Folk som sitter ute i en park på en sten.
Två kvinnor pratar med varandra på en gata.
En ung kvinna som har ett genombrott på en stor mur.
Två tonårspojkar tävlar, den med långt hår vinner.
En man som bär en grön långärmad skjorta springer.
Ung pojke i vit skjorta kör på ett spår som håller en markör.
Flera personer står vid en busshållplats.
En livlig stadsscen med många olika typer av fordon antingen parkerade, eller flytta längs på motorvägen.
Ett barn i grön skjorta cyklar.
Två hundar jagar varandra i gräset
En man bär en väldigt konstig hatt.
Ett actionskott av en unge i grönt utför ett skateboard trick från några steg.
En grön cykel står parkerad bredvid en dörr.
En kvinna med svart hår med en ärmlös klänning står bredvid en bil.
En flicka sitter på en smal kanot.
Damen med mörka nyanser på är i ett samtal med sina vänner.
Man i blå skjorta och röda shorts står på trottoaren.
Många rosa och lila ballonger trängs in i ett utomhusområde som en kvinna med ett paraply går förbi.
En skara människor i ett gathörn, tre pojkar med sina skjortor instoppade.
Människor befinner sig i ett område där belysningen lyser upp området.
Folk går på en gata på natten.
Två män och en kvinna promenerar längs gatan förbi varuhusen.
Det här är en man som skyfflar snö, bredvid en bil.
Ett ungt par som går ut vid en vägg med graffiti på och en ljusblå äldre modellbil.
En ung man med retro frisyr väntar bredvid en bil.
En grå och brun hund hoppar från en brygga in i en sjö
En man tar ett foto av en kvinna som bär en orientalisk hatt på en liten docka.
En pojke med en vit skjorta upprullad visar sin mage och ler.
En man i hatt sitter i en stol.
Ett par tar sin egen bild framför Arc De Triomphe, från andra sidan gatan.
En stad på natten med människor som går runt.
Man med ryggsäck på promenader ner för en gata, röd informationsstånd i bakgrunden.
Ett par går nerför en gågata på natten.
Gult ljus badar flera restauranger som sitter utanför en liten fransk restaurang.
En kvinna på en offentlig marknad skär en kyckling i små bitar
En man tittar på saker till salu på gatan.
En grupp människor samlas på ett köpcentrum.
En kvinna i baddräkt sitter på en brygga över en vattenförekomst.
En grupp människor står på trappan framför en byggnad.
En skara människor väntar på toppen av trappan utanför en byggnad.
En kvinna i batmanskjorta går nerför strandpromenaden.
En massa människor med fokus på en kvinna med långt blont hår och en svart skjorta.
Flera människor köper mat på en asiatisk matmarknad.
Motorcyklist racing på ett spår med en gul smuts cykel och en Kawasaki-märkt grön annonsskylt.
En man med stor mustasch och lila hatt.
En hona går uppför en trappa med vatten till vänster.
En flicka håller i en kamera och gör en handgester.
Två personer kan ses på avstånd i en gränd mellan två stora byggnader.
Dam i vit skjorta med en grön väska poserar för kameran
En äldre kvinna klädd i rosa går och håller i en tidning.
En tjej med vit klänning poserar för kameran.
Ett äldre par poserar med en motorskoter, medans de bär renässansfestivalkläder.
Mannen funderar över sin situation under en promenad genom gården.
Ett antal personer går över framför en rulltrappa.
En snowboardåkare i luften, med en färgglad dekorerad bräda.
En man utan skjorta som sitter på en stol på en flodbank och pratar på en mobiltelefon.
En körgrupp reagerar på skott som avfyrats under en ceremoni.
En asiatisk man i korta shorts och knäskydd joggar nerför gatan.
En motorcykelförare gör en skarp sväng.
En man i en hatt med en kamera och en dam med en skylt.
En man som bär en fängelseoverall är att få sin bild tagen
Äldre man i vit skjorta och svart slips klädd i svart basker och går nerför gatan.
Två kvinnor delar paraply på trottoaren.
Två pojkar på skateboard framför en staty av en soldat på en häst.
En snowboardåkare gör ett hopp i en tävling.
En cyklist med långt blont hår som äter en glasskon.
En kvinna i blått pratar med en fruktförsäljare på gatan.
En grupp snowboardåkare flyger över en kulles krön.
Två kvinnor, en rosa klädd och en orange klädd i kökssysslor.
Ett ungt par håller hand när de går längs en stadsgata.
En man och kvinna njuter av utsikten över staden.
Ung kvinna med scrabble skor och vita fälgade solglasögon pratar och ler på mobiltelefon medan du öppnar paketet.
En man i vit skjorta röker medan han ger instruktioner.
En ung pojke som äter en liten kaka ligger i en kundvagn fylld med matvaror.
En man i svart skjorta är under en eldklot.
Tjejen med den rosa träningsutrustningen gör en flip.
Folk använder crosswalk på storstadsgatan.
En liten flicka sparkar en boll framför ett fotbollsnät.
Kvinnan tittar noga på skor hon gillar.
En ung man och kvinna går på en trottoar bredvid en vit byggnad.
En man som sitter ensam på ett picknickbord framför en gul lastbil och äter lunch.
En familj, dotter i mitten, går nerför gatan.
En man och hans son går förbi en vuxen videobutik.
En äldre man med grått hår står utanför en affär.
Ett barn i röd skjorta sitter på sin fars axlar.
En ung blond kvinna går genom en gata med en svart handväska.
En ung flicka håller ett basebollträ över axeln
En knubbig man rider iväg nerför gatan på en cykel.
Män och kvinnor i en militärparad.
En grupp människor i orange kostymer står runt stora paket.
En pojke sitter på gräset nära en geometrisk skulptur.
En person på en mobiltelefon står vid ett fönster i ett högt tak rum med svart vitt en röd bricka.
Folk är på en avsats utanför en byggnad.
En tonåring utvecklar sin skateboardteknik framför en vacker, utsmyckad byggnad.
Två personer kysser varandra på gatan i en väl upplyst stad.
En kvinna som sitter på trottoaren får ett armband som ges till henne av en annan kvinna.
Den här damen bär en rosa skjorta och tutar sin gitarr
En stor grupp cyklister rider nerför en gata.
Sju brandmän tittar upp mot en byggnad.
En polis är på väg ut från ett område med polisband medan åskådare tittar.
En grupp människor står på en trottoar.
En man med glasögon läser genom en meny på en restaurangs uteplats vid sjön.
En man med ett vapen som ligger mot en vägg.
En munk i en gräddtunika som står på en marknadsplats.
En gammal man med en käpp som står utanför.
Sex personer sitter vid fönstret i en restaurang och gör sig redo att beställa.
En manlig figur som står och kikar över en vattensamling.
En man bär en rutig hatt, en klocka, jeans, många tillbehör, och en skjorta med en vit cirkel och nummer fyra i mitten.
En grupp människor tittar bort från ett observationsdäck.
Två män som talar medan de tittar över räckena över en flod.
En man tar en paus från sin vandringsresa.
En man går på en trottoar framför en byggnad.
En ung blond dam tar en cigarett medan hon går.
En man och en kvinna bär hjälm medan de kysser varandra på gatan.
Ett gammalt par går nerför gatan och håller varandra i handen.
En flicka i rosa jacka går först nerför en röd rutschkana.
En man i jeans och sandaler som ritar i en vägg.
En man i vit T-shirt och blå overall går nerför gatan.
En äldre man som gick förbi en byggnad täckt av graffiti.
En vacker stad skjuten med en fontän och en dam sitter på några steg.
En man sitter på ett fartyg och läser en tidning.
Det är en kille som barbecuing och han bär glasögon och en röd hatt.
Det här är en ung pojke på en strand som håller i en pinne.
En ung flicka kör en rosa leksak Cadillac bil.
Många människor tittar på en man i gult gör djurballonger.
En familj på tre avkopplande mitt på dagen.
Mannen på trottoaren sitter på en motorcykel.
En kines knuffar en rullstol utan någon i den på en hektisk kinesisk gata.
En tjej med varma rosa tånaglar och baddräkt ligger på en varm rosa handduk.
En kvinna i en blå bikini övredel går.
En flicka tittar på sportspelare av en vägg täckt av graffiti.
Tre män sitter på trottoarkanten framför en närbutik.
Två män sitter på trappan utanför.
En brud och en man ses utanför byggnaden när de har gift sig.
Ett par i affärskläder sitter på ett hörncafé med al fresco middag.
En familj sitter i en vinterträdgård med trädgårdsstolar och har picknick.
Gamlingen står med vit t-shirt och hatt.
En man tar tag i stöd när han går på en ställning.
Leverantörer serverar mat på gatan.
En kvinna i vit hatt och en röd och vit randig skjorta som sitter på en vägg.
En asiatisk kvinna i vit skjorta som sitter i en blå stol.
En person som målar en väggmålning på sidan av en byggnad medan människor står och tittar.
En publik väntar på att interagera med en del människor på en inomhusplats.
Ett fattigt bostadsområde med en kvinna i svart med vit huvudbonad på avstånd.
Två män står utanför bredvid en byggnad.
Tre poliser står runt någon i en grå tröja med ränder.
En man med hatt som lutar sig mot ett inlägg och läser en tidning.
En man som sitter och en kvinna som ligger i hans knä kysser varandra.
Fyra personer i fallskärmshoppning i ett plan högt över jorden.
Två kvinnor bär bikini toppar och mycket korta shorts medan de går nerför gatan.
Det är mörkt ute och två kvinnor står här.
En grupp människor går i en avslappnad linje över en stenlagd innergård.
Tjej med polotröja och kille med stor buskig frisyr väntar på att korsa vägen.
En ung man i en randig hoodie tittar på en konstnärlig Levi annons som säger "Vi är alla arbetare."
En asiatisk flicka som står utanför en byggnad.
En kvinna sitter i hörnet och äter en smörgås.
Människor i traditionell militärtjänst och två människor ridande elefanter någonstans i Sydostasien.
Två män kliver sida vid sida på trottoaren längs en röd målad vägg.
Skolbarn klädda i gult.
En kvinna i svart, sedd bakifrån, sitter bredvid en vattensamling.
En blond kvinna som sitter med benen korsade med slutna ögon.
En man med svarta byxor och hatt sover på en bänk framför en historia byggnad.
En grupp män som står ovanpå en ubåt
En grupp människor som är klädda snyggt slappnar av tillsammans på grönt gräs.
En liten pojke med gröna och röda kläder och sandaler, som hukar sig ner på en trottoar.
Två män som bär röda byxor och håller fast vid en vertikal stege, verkar göra akrobater utanför en byggnad.
En ung dam sitter nära hem med solpaneler.
En blond tjej med blå rock sätter på hjälmen för att cykla.
En väggmålning med ögon och händer säger "stoppa våldet, vi hjärta en säker NY."
En garvad kvinna cyklar medan hon bär en vit bikini.
En turistbåt på en flod vid en falsk gammal byggnad.
En kvinna sitter på en moped i en affär.
Tre personer står på en brandstege.
Två personer klädda i idrottskläder går nerför gatan, medan den längre av de två håller en basketboll.
Två unga män som pratar framför ett basketbord i Penn State.
En man lutar sig över en bil med skägg som tittar på kameran medan han arbetar på en bil.
En kvinna med rött hår som tittar åt vänster.
En man i en blå tröja och svarta byxor lämnar en nyhet och livsmedelsbutik.
En mamma som knuffar en barnvagn och håller handen på ett litet barn.
Brun hund med öppen mun stående mitt i grönskan.
En grupp människor slappnar av vid några bord.
En man i baseballmössa och solglasögon står i en godiskiosk.
Fem personer står under en asiatisk valvväg.
En grupp människor samlas och tar bilder i en innerstad gemensam mark.
2 Kinesiska människor bär traditionella kläder
Tre män i hårda hattar, ett par och ett barn ser ner på något.
En man sitter på stranden bredvid en stolpe.
Ledande sångare i ett band har ett papper och en mikrofonstativ med detta band som spelar bakom.
En kvinna med shorts och höga klackar lyssnar på något på sin telefon.
Flera människor sjunger till mikrofoner och dricker.
En fri löpare hoppar en rail.
En man, i en blå jacka, sitter i regnet under ett grönt paraply.
En lång stadsgata omgiven av stora byggnader
En utsikt över folk som går på gatan nedanför.
En kvinna som hular i en röd skjorta.
En man utan tröja står bredvid en container utanför.
En grupp barn som leker med rekvisita
En ung hockeyspelare som spelar i isbanan
En kvinna undersöker ett prov genom glasögonen på ett mikroskop.
Ett par lägger armarna runt varandra och går längs en lång korridor som stöds av stenpelare.
Ett barn i riddarkostym som blir fotograferat.
Två personer omfamnar framför en byggnad med logotyp på byggnaden som säger Monk Kok.
Det är en våg på väg att ta ner en surfare.
En man i en bollkeps står på en korsning med en flagga i en fullsatt stad.
En kvinna som uppträder på scenen med en mikrofon.
En man går nerför gatan framför en vit skåpbil.
Två motståndare spelar på en plan.
En person som flyger en hängglidare över en stad.
Folk filmar en kvinna som rapporterar.
En man i en kanot kastar ut ett fiskenät i vattnet.
4 personer verkar flytta olika föremål från en byggnad
Män och kvinnor går längs en trottoar bredvid en trädgård.
En ung pojke står i en knapp-down skjorta och shorts.
En flicka fotograferar på en fin gräsmatta medan andra sitter bredvid henne.
Tre unga män möter en äldre man med visselpipa.
En äldre kvinna i blått och rött korsar gatan i en korsning.
En pil som pekar på en man i en vit hatt som går förbi.
En kvinna går med sin cykel bakom två personer bär paraplyer.
En flintskallig man som går bland pelare på en trottoar.
Det finns människor som går på en hektisk nattgata med skyltar som lyser vägen.
Tre unga barn som sitter vid en vacker utsikt.
En grupp män och kvinnor som hänger på en klippa och spelar in landskap.
Person i en grön huva tröja, tittar på utsikten.
En stor grupp små barn står på rad, medan flera vuxna tittar på.
En person sitter framför en graffititäckt vägg.
En grupp små skolpojkar som bär uniform tar en paus framför en stor apstaty bredvid havet.
Folket korsar gatan mot en restaurang.
Två svarta och vita hundar på sandstranden slåss om en lång pinne
Två små pojkar lagar en liten cykel.
En jockey rider en brun häst på en trottoar vid en vattensamling.
En busshållplats innehåller många personer med intressanta föremål.
Grupper av människor går nerför en smal gata, en kvinna som bär en svart skjorta bär ett vitt paraply.
En man i en skjorta som läser Hippie Killer ler mot sin flickvän i en Return of the Living Dead-tröja.
Några personer går i ett vattenområde.
Den här mannen tänjer på sin halsduk och jublar.
En ung man går genom en pöl utanför med en blå trehjuling cykel står parkerad i samma pöl.
En man som står nära en pinnestruktur.
Dessa små flickor är i kinesiska geisha kläder och smink, håller röda paraplyer.
En skjortlös liten pojke skyddar sig lekfullt från en brandmotors sprej med ett paraply.
En man i idrottskläder som böjer sig ner för att binda sin sko.
Grupp av människor på däck av strandhus
En kvinna i röd skjorta som står på en öppen gård och tränar med en man i vit skjorta och byxor.
3 personer rider motorcyklar nerför gatan.
En man med en mask med gröna dreadlock och blå handskar står framför en kvinna i en brun kofta.
Tre cowboys på hästar arbetar tillsammans för att repa en kalv.
Den stora vita kon är dekorerad med en röd trådkula.
En tonåring i röd skjorta cyklar.
En kvinna med stora leopardörhängen tar en video.
En kvinna poserar med en skråma på ett torg.
Ett barn jagar ett annat barn som håller i en fotboll.
En kvinna i röd skjorta och hatt röker under ett religiöst märke.
Två hundar brottas över en bit svart material.
Många protesterar när de går nerför gatan.
En ung pojke i gröna byxor står ensam på en väg.
En kvinna sitter vid vattnet nära två elever.
En dam med blått hår sitter och spelar gitarr framför en blå vägg.
En kvinna i randig skjorta pekar på något med sitt blå paraply.
En stadsgata där en kvinna med brun väska och vita kläder passerar en utställningsbutik.
En karikatyrkonstnär sitter under ett rött och vitt randigt paraply.
En ung blondhårig pojke med ett nummer på framsidan lutar sig mot ett räcke.
En kille på en motorcykel i en gatubelysning.
En grupp av tre asiater som står mitt i en storstad och diskuterar något.
Ett uppspelt barn som springer i ett lopp.
Stadens trottoar med affischer på en vägg, flera människor går förbi med stadsbyggnader i bakgrunden.
En man i svart skjorta skålar en orange bowlingboll.
En man lutar sig framåt på ena foten i en bowlinghall strax efter att ha släppt bowlingbollen ur handen.
En kvinna i brun skjorta som sitter på en bänk.
Ett par går upp för trapporna till en bro i en innerstad av en stad.
Brunettkvinnan sitter på en stol i hörnet av gatan och läser.
Fyra personer sitter utomhus vid ett vitt fyrkantigt bord när en man i en randig rosa skjorta står och pratar med dem.
En ung man med glasögon ser frustrerad ut i en tvättomat.
En flicka väntar på att gå över gatan medan hon tröstar ett barn i en barnvagn.
En kvinna går längs trottoaren framför en spegel
Ett barn och en vuxen går längs trottoaren.
Två personer sitter framför en dator medan de bär solglasögon.
En man rider en wakeboard fastsatt i en fallskärm.
En ung man i svart t-shirt med en grön hatt stående.
Två kvinnor i baddräkter vid en bänk stirrar upp på en gigantisk vit ballong.
Fyra män går nerför gatan i sin orange klädsel.
En ung man är skysurfing med en bräda som har målat en orange flamma skalle
En man parakiterar på en vattenförekomst.
En kvinna som bär en mörk topp och mörka solglasögon går i kilklackar och gör ett ansikte.
En man som kör maraton pratar med sin vän.
En man i vit t-shirt sitter på motorhuven på en bil.
En kvinna knäböjer på marken och tar ett fotografi.
Gamla kvinnor som använder en vandrare för att gå ner för trottoaren.
Den äldre damen i den vita kjolen bär rosa skor.
En skara människor som kommer nerför trappan från hovhuset.
En liten pojke som somnar i sin pappas knä på en grön gräsmatta.
En blond kvinna med 40-tals frisyr och leopardtryckt skjorta.
En man och en kvinna går över gatan klädda i formella kläder.
Protester är i bakgrunden av detta foto medan en tidningsvisning är i förgrunden.
Folk går nerför gatan, par i förgrunden med paraply.
En flicka i klänning går nerför gatan och gatan är full av träd.
En parkeringsplats i staden med folk som går genom den.
På äldre asiatisk man i en gul knapp ner tittar på kameran.
Svart man jonglera en basketboll, bowlingboll och en tennisracket.
Arbetaren bär en mask för att skydda ansiktet mot kryddiga chiliångor.
En kvinna håller upp kjolen på sin klänning.
Två gatumänniskor och en hund som sitter på marken och en håller en "oturlig" skylt.
Folk samlas på en gata.
En gammal man sover på gräset vid foten av ett stort träd.
Två arbetare med hattar står på ett fält.
Asiatiskt par med två barn tittar på frukt och grönsaker i en monter.
En man i mörka kläder sitter på en bänk framför en lastbil.
Två män klädda i vita dräkter och röda capes rider cyklar medan de bär stavar toppade med skallar.
Några personer står nära vita pelare framför en gul vägg.
Två män målar modern väggmålning på en vägg med en inrullande gångväg.
En man med tatueringar med skateboard ger tummen upp på trottoaren.
Kvinnor klädda i röda och svarta klänningar går i en cirkel framför en butik som en liten publik tittar på.
En man i gul t-shirt har en stor videokamera.
Flera indiska kvinnor i färgstarka kläder arbetar.
En grupp människor har ett samtal utanför en byggnad.
En del människor samlas framför en byggnad med affischer upphängda på väggarna.
En lockigt hårig man spelar gitarr vid en ceremoni medan folk tittar på.
En Cola lastbil kör förbi en blå lastbil parkerad på sidan av vägen.
En kvinna som går med matvaror och går förbi graffiti
En flicka klädd i svart med en handväska på armen ler mot en man i ett rum med massor av desserter på bordet.
En man med vit skjorta och svarta shorts går förbi några gamla byggnader.
En man i vit skjorta och en kvinna i orange topp sitter tillsammans på stranden.
En man väljer en tomat på en marknad.
En man är i luften och utför ett trick på sin cykel mot en molnig blå himmel.
En man i blått tar sig genom en folkmassa under ett lopp.
En man som bär rött sitter upp i luften på en plattform.
En flicka som sitter på en sten och tittar över sjön.
En man går nerför trottoaren till sin destination när han når in i fickan.
En cowboy som kastas av en häst på en rodeo.
Smickrande barn med fåniga blå hattar på huvudet.
En grupp kvinnor klädda i lila samlas nära en lastbil.
Flickan bär lila kläder och svänger upp och ner.
En man som pumpar bensin på sin mobil.
Tre hundar leker tillsammans på det gröna gräset.
Tre springande män deltar i ett maraton.
En kvinna i grön skjorta kör ett lopp och tittar på sin klocka.
Folk går nerför en pub-laden gata omgiven av affischtavlor.
En man går längs en kullerstensstig, bredvid en stor blå vägg.
Kunderna väntar på att få lite mat.
En man som bär shorts och svarta skor uppträder framför en publik.
En grupp människor tittar på sandskulpturer.
Någon som ligger på en stor solbränd soffa utanför bredvid en parkeringsmätare
En man pratar på sin mobil i enrum.
En hona i en blommig skjorta med en brun meny.
Kalifornien springer tillbaka och tar hand om det.
En sömmerska arbetar för att passa modell skyltdockor i hennes mörknade studio.
Kvinna bär färgglada halsduk bland människor glatt flin.
En brunhårig kvinna med röd skjorta, en blå ryggsäck och solglasögon på huvudet.
Brunett kvinna i en vit skjorta, stående framför en disk.
En asiatisk man förbereder sina produkter i sin monter för den dagliga marknaden.
En kvinna med tunt hår arbetar i en köttbearbetningsanläggning.
En person som slår en boll i en omgång Cricket.
Två flickor som går under ett lila paraply.
En kvinna med en stor handväska som vilar sin fot mot en vägg.
En man målar en livlig orange och gul vägg.
Två manliga idrottare i svarta skjortor springer längs en gata.
En yong kvinna i grå skjorta har ett halsband hon har på sig.
Folk klädda i formella kläder förberedda för en händelse.
Vissa deltar i en road race.
En svart hund och en vit hund leker med varandra och en grön boll.
Ett litet barn klädd i en vit dräkt.
Någon som inte bryr sig om jorden var här.
En äldre kvinna i klänning står nära buskarna.
En person sitter i en park medan han spelar ett litet instrument.
En skara människor som går genom en promenadväg av olika slag.
En ung man står utomhus framför elektronisk utrustning med armarna ihopfällda medan en annan man i bakgrunden bär hörlurar.
Många människor går längs en fullsatt gata.
En dam knuffar en barnvagn medan en man bär ett barn på axlarna medan han går och bär Labor Day 2010 blå t-shirts.
En clown delar ut amerikanska flaggor och underhåller några barn.
En ung blond pojke som rider en röd, vit, blå och gul cykel med amerikanska flaggor på.
En man och en kvinna med ryggsäckar är utanför.
Folk går ombord på ett blått, vitt och guldtåg.
Två mörkhåriga unga kvinnor klädda i t-shirts springer i ett lopp.
En svart hund jagas av två bruna hundar på stranden.
En kvinna som pratar med en person utklädd till frihetens staty.
Ett barn sitter på en motorcykel som som en amerikansk flagga kommer ut bakvägen.
En hånad frihetsstaty står i folkmassan.
En kvinna i röd skjorta vinkar medan hon står bakom en annan kvinna med svart hår.
En äldre man sitter i en stol i en gränd.
En man som gör fönstershopping för sina skor i en sportaffär belägen i staden av vinklar
En man bredvid en häst sitter i en stol och säljer konstverk.
En brandman i Seattle står framför sin lastbil.
En brandman ser sig omkring i djupa tankar.
Två brandmän med "Seattle Fire" på baksidan av sin utrustning möter sin lastbil.
Två män springer i ett lopp, sida vid sida.
Utanför ett företag visas med en soptunna och fyra personer går runt.
En dykare spelar trummor.
En man som sitter vid ett fruktstånd pratar med en pojke i en bokpåse.
Leverantörer säljer frukt på en utomhusmarknad under ett olivträd.
Två brandmän gör sig redo för en brandbil.
En brandman klädd i växel ser förbryllad.
En grupp mörkklädda män samlas utanför och talar entusiastiskt.
Många i vita skjortor går nerför en gata.
En kvinna som bär röd skjorta sitter bredvid andra på en trottoar och håller i en kamera.
Två unga män i kamouflageställning i gräset.
Vad är en resa till parken utan att besöka snackbaren?
Två flickor uppfostrar en annan flicka i luften.
En kvinna, som bär en färgglad bikini, vilar bredvid det blå vattnet.
Ett par sitter utanför en anläggning.
En asiatisk kvinna i röd polotröja tittar över en disk.
En man som går nerför en skuggig gata med en shoppingväska.
Hon solar sig med sitt lilla gula paraply, när hon visar upp sin fina långa klänning.
Landsmusikgruppen - Sugarland, framförande.
En äldre person som vaknar ute på dagen med solglasögon på.
En kvinna i vit klänning med blå smycken håller i en tupp.
En man i vit skjorta, på en skoter väntar på trafik.
En man bär handskar och en hjälm.
En man som sitter framför en vägg av graffiti.
En hårt arbetande man talar sitt sinne in i sin megafon.
Tre personer i en liten båt bredvid en träbrygga där två andra människor står.
En tjej i ljusa kläder som dansar med en hulahoop.
En kvinna som bär en rosa, prickig ryggsäck håller ett litet barn.
Fyra kvinnor går genom ett konstgalleri.
En kvinna med orange skjorta går förbi en 1 timmes fotobutik.
En äldre kvinna staplar tallrikar att placera i sin vagn.
Vit man med långt grått skägg, bär svart hatt och lång svart kostym när han går nerför gatan.
På en nöjespark eller basketplan.
En man i den blå skjortan tar ett foto med en familj han träffade på semestern.
En kvinna och en grupp barn som lever i fattigdom.
En liten pojke med randig skjorta som går genom gräset nära några träd.
En pojke svänger på en pinata under en utomhus familjefest.
Smickrande barn sitter på betongplattan och visar ett litet föremål i sina händer.
En man i grå skjorta håller i en hammare.
En kvinna i svart lutar sig över en flerfärgad bänk medan hon tittar in i en röd hink.
Tre kvinnor rider i en vagn.
En ung kvinna söker igenom sin väska nära ingången.
En tjej som bär solglasögon och en orange tank topp hula hoops.
En kille går med eld i handen och en CGT jacka på när två killar tar hans bild.
Män som bär röda skyddsvästar och bär skyltar går nerför en gata där en explosion har inträffat.
En grupp kvinnor, några med hijabs, samlas runt en kvinna som sitter på en moped.
En gammal kvinna som står nära påsar med saker.
En kvinna med fjädrar i håret och en hennatatuering i ansiktet tittar utanför skärmen.
En man, kvinna, ett barn som sitter på bänkar och väntar på bussen.
En kvinna som håller i en svart väska håller fast vid ett stängsel.
En flicka ler utanför en affär.
En man i mörkblå skjorta och röd ryggsäck går vid en graffititäckt vägg.
Två män står på trä, båda bär hattar.
En kvinna med en shoppingväska som går mot en gata.
Lunch utomhus en solig dag.
En kvinna i jeans och en blå skjorta står utanför och röker en cigarett.
Kvinnor går nerför gatan i jeans, svarta högklackade stövlar och en beige handväska.
Det finns grönsaker till salu på en marknadsplats och en man trycker ner sin lastade cykel.
En kvinna och en man dansar offentligt
En brunett i en orange skjorta som leker med en grön och vit hulahoop.
En man som går med ett protesttecken.
En parad äger rum och människor är klädda med ljusa färger.
En flinande man med spikar av flerfärgat hår och stora öron-piercing
En asiatisk man studerar insidan av en glasbyggnad från gatan.
En flicka skriker när hon kommer från vattenrutschbanan.
En man och en kvinna kysser varandra i hörnet av en gata.
En man går längs trottoaren med en ryggsäck och ett paket.
En man ser uttråkad ut medan en annan man tittar genom två juvelerarmikroskop medan ett barn är underhållet.
En halvnaken skyltdocka är poserad i fönstret.
Fem personer med dykutrustning samlas i lugna vatten.
En kvinna böjer sig över för att titta i sin väska.
En kvinna i leggings och tunika, läser en flygare på en ljusstolpe.
Par delar mellanmål på offentliga monument på solig dag.
En liten grupp hundar drar en vagn full av barn som är täckta av blommor.
En pojke i en blomstervagn dragen av hundar.
En kvinna och hennes dotter väntar på sin skjuts efter att ha fått mat när två personer går förbi dem.
En kvinna går förbi en fontän med palmer i bakgrunden.
Tre personer sitter och tittar över ett dräneringsdike bredvid en krokodilvarning.
En kvinna i vita byxor som håller ett barn tittar på havet.
En ung kvinna klädd i grönt och brunt sitter på trappan med ett papper i knät.
Person fallskärm, med solen och himlen i bakgrunden.
En kvinna som står bredvid sin cykel och väntar på att få gå över gatan.
En man kör ett mycket litet fordon.
En man i en beige och vit randig skjorta, bruna shorts och skor med en hand på ansiktet och en fot upp ser framåt.
Folk sitter och går längs gatan i en stad.
Två kvinnor sitter i baksätet på en lastbil och äter.
En man tar sin katt på en promenad i stan.
Tre solbrända män på sidan av ett berg tar en paus från att gräva.
Två personer lounge i ett stort utomhusområde.
En äldre kvinna med en väska som går under en flygplatsskylt.
Två personer står framför en byggnad med graffiti som lyder "Boss Life".
En kvinna står vid en cykel, framför en affär och tunnel.
En polis skriver en biljett för dålig parkering.
En flicka som sitter vid ett skrivbord i ett bibliotek lägger sitt huvud på en bok.
Två män spelar trummor framför en folkmassa.
Många ungdomar sitter på en vägg och hänger tillsammans.
En kvinna med vit blus går bort från en byggnad.
En grupp surfare paddlar ut i vattnet.
Man med rött hår i gröna byxor under ett paraply poserar för en bild.
Två pojkar leker på en stad gata; den med glasögon ger en V-signal till kameran.
En kvinna sitter på konkreta steg bredvid en teckning av ett hjärta.
En man i blå skjorta och svarta byxor promenerar förbi en irländsk pub.
En man sitter på en blå skoter på gatan.
En kvinna sminkar sig själv.
Ett barn med blont hår står nära sin cykel på en osökt väg.
En man lutar sig över för att kyssa en kvinna på en cykel nära en palm.
En hund ser ut över grönt gräs och blommor.
En grupp mestadels yngre personer som hänger i en bubbelpool på hotellet.
Byggutrustning framför en byggnad med en väggmålning av en man som lyfts av svarta fåglar.
En dam cyklar på ett trädäck vid stranden.
En man som sitter med sin lilla hund.
Fyra hanar i olika åldrar täljer ut mönster på stora vita plattor i en rörig, öppen för luft verkstad.
Röken kommer från ett jetplan i himlen.
Två män med stegar arbetar på ett staket.
En ung backpacker sitter på en bro med utsikt över en flod.
En grupp människor fotograferar samtidigt något uppåt.
Arbetare bär sina hattar på en avsats.
Tre blondiner klädda i svartvitt går över en bro på dagen.
En grå bil väntar på att ljuset ska bli grönt vid en korsning.
En man som bär en grå hjälm bredvid sin moped i ett hektiskt område.
Två afrikanska soldater går in i en stor stenbåge, en man som ger tummen upp.
Män i armén som håller i vapen.
En man med blå blazer går ut.
En ung pojke tittar på kameran medan han bär en New York-hatt och en svart och vit randig skjorta.
En pojke på en grön cykel får ett samtal.
En kvinna i grå klänning poserar utanför Louvren.
En gatuscen av människor på scooters.
Ett barn i vit skjorta kommer ut ur en sving i luften.
Två honor omfamnar varandra.
En person i laxfärgad skjorta tar en bild av något ovanför dem.
En kvinna som tittar upp på en fullsatt gata.
En man som bär en blå tröja och en solbränd strumphatt röker en cigarett.
En man på en cykel går en hund längs en strandpromenad.
En dam i blå skjorta som gör ett lustigt ansikte på en liten flicka som biter något i en restaurang.
Ett par går förbi ett café där ett annat par sitter utanför.
Två gatuförsäljare sitter på trottoaren och väntar på kunderna.
Tjejen manövrerar en cykel genom en tältsats utanför.
En kvinna som bär vit träningsoverall sträcker foten över huvudet.
En clown håller öronen med en ballong i vänster hand.
En gammal man pratar med en annan man som bär militärdräkt och är nära en apa.
En man som cyklade med tidningar i korgen.
En ung pojke tittar tillbaka på kameran medan han sitter på en röd skoter.
En elev rusar till lektionen samtidigt som han har hörlurar på sig.
En dam i rosa kappa som går med ett litet rosa paraply i handen.
En professionell fotbollsspelare försöker korsa bollen, medan en annan försöker göra tacklingen.
Två kvinnor står runt ett täckt bord utanför omgivet av vackra blommor.
En kvinna i en svart mössa tittar upp på en skäggig man.
En man som står på gatan och njuter av arkitekturen i en byggnad.
En kvinna poserar utomhus med ett designparasoll.
En grupp asiatiska kvinnor klädda i färgglada kläder och håller fans.
Åskådare observerar som London Arsenal FC utövar fotboll på deras plan.
En liten person håller en gul flagga med en röd logotyp på sig.
En man i orange pratar på sin mobil.
Kvinnan i rosa och grön tank topp lyssnar på en man i grönt bär en blå ryggsäck.
Flera människor är sysslolösa runt en plaza i skuggan.
En äldre skäggig vit man med blå skjorta och röd jacka tittar ner på en korv han håller.
Två gamla män i polotröjor.
En man i vit skjorta och byxor håller i ett rep och tittar upp.
Det är en parad med folk klädda i kostymer.
En man som bär en grön skjorta och bär en shoppingväska läser tidningen i ett stadshörn medan en kvinna tittar på.
Folk går över en korsning.
En gammal man i en vit tank topp kliar huvudet.
En medelålders man hukar sig i ett smutsigt rum.
En man med paraply står på en bergssluttning och det regnar.
Ett barn som bär hatt och ryggsäck går genom stan.
Många manliga arbetare står utanför en byggnad i gröna och blå kostymer.
En kvinna i en svart tank topp hula hovar.
En man går nerför gatan bredvid en vägg med en stor mun målad på den.
Kvinnan med scarfen tittar på när mannen lagar mat.
Två män bakom disken i en söt affär medan två människor tittar på godis.
En kvinna använder en sked för att servera mat.
Ett ungt par blickar in i varandras ögon medan de rider på en rulltrappa i en shoppingvagn.
En man i svart skjorta går sin hund under solnedgången.
En man kollar sin telefon när han går sin hund längs piren.
Liten medelöstra barn i typ av trä underjordisk grotta.
Ett litet asiatiskt barn rider på baksidan av en kvinna som bär hatt.
En sportbar där du kan titta på spelen.
Ett asiatiskt par sitter på en träbänk i ett skogsområde och läser och ser sig omkring.
En flicka och ett litet barn tittar åt olika håll på en trottoar.
En gatuförsäljare klädd i kockhatt och flera människor samlades runt honom och hans vagn.
Två kvinnor i rockar tittar på en utomhus smycken display.
Två män är på en strand och tittar på avstånd.
Mannen i den blå jackan gick förbi telefonkiosken.
En kvinna i skjorta korsar gatan en molnig dag.
Två män går på stranden med gitarr i handen.
En man i en ljusgrå t-shirt kör en ljusröd Coca Cola lastbil.
Två män och två unga kvinnor jobbar på en blå cykel.
En fotograf står i skuggorna framför en vägg täckt med graffiti.
Folk tittar på föremål på en utomhus försäljning.
En kvinna i orange skjorta och vita byxor går i kyrkan.
Barn vilar och går uppför många trappsteg.
En vithårig man och en brunhårig kvinna går tillsammans och håller varandra i handen.
En servitör står vid ett bord.
Två personer står framför ett matbord.
En man som står med sina ögon nedslagen.
En asiatisk man som hukar sig på gatan med tillhörigheter.
En kvinna som njuter av en drink i solen.
En person cyklar i en tunnel.
Vit hund vid vattenbrynet.
En man i vit skjorta äter, står bredvid ett staket.
En man böjer sig ner på en sten.
Fyra män, i röda hattar och orange uniformer, går nära en häck.
Två män spelar instrument på gatan för att underhålla förbipasserande.
En man väntar vid tunnelbanestationen på att tunnelbanan ska anlända.
En äldre man i kostym låser sin cykel.
En gata med en ensam man i mitten.
Hunden stirrar på något med en leksak i munnen.
En man klädd i svart och vitt står på sidan av gatan och äter en glasstrut.
En man på en fruktmarknad som tar tag i lite frukt.
Studenter som har rast efter att ha tagit ingenjörsexamen i sin skolsal
Två män i kostym och hatt går tillsammans.
Fotgängare samlas i ett gathörn, framför Lyppens och Schipper butiksfront.
En liten pojke i gul t-shirt lär sig att skriva.
Den mycket trötta svarta damen bar sin nya röda blus, när hon red hem på bussen.
En grupp människor samlades och tittade på två män som lyfte en kvinna på en träsåg.
En ung kvinna tycks dras ut ur en dräneringskanal av en stol som är fäst vid en trä 4 av 4.
En person lyfts upp ur vattnet med en gammal lyftare.
En grupp på tre äldre och tre yngre personer står samlade i en vattenförekomst.
Två flickor i en blomstersäng med armarna utsträckta.
En kvinna är i luften medan hon vaknar av en våg.
En man läser en tidning medan han väntar på ett tåg.
Tre personer sitter och tittar ut på vägen och håller en karta mellan dem.
En man utan tröja på knyter en gul genomskinlig väska stängd.
Tre vita män klädda i tillfälliga kläder, en i blå overaller, en i orange bollmössa och en i gul skjorta går över en gul ställning.
Asiatisk kvinna i publiken, bär svart väska med "smärta" och spetsade knoggrafik.
Två små flickor bär ljusa klänningar blåser bubblor med bubbelstavar.
En man och en kvinna, båda klädda i svart, dansade tillsammans
Kvinnlig målare målar på en vas med tre personer som tittar på henne.
En man med en brun halsduk som blåser rök.
En förvrängd bild av en ung pojke som springer
En asiatisk tjej som äter en korv på ett matställe.
Två personer, en i lätta jeans och en randig skjorta, spelar pool.
En flicka städar trägolvet med en swiffer.
Fotbollsspelare klädda i röda och vita uniformer går på ett fält.
En man som satt fast i trädet.
En stor klass av utexaminerade som bär dräkter och murbruksbrädor väntar på sina diplom.
En man som tar en bild från en bås med linslocket på.
Tre män i shorts står på parkeringen i en byggnad märkt en "fabrik".
En hand håller en utsmyckad metallbit.
En ung pojke i jeans och en blå skjorta bär en blå hjälm.
En ung kvinna rider i en bil.
En man sitter och funderar på något medan en man sitter över sin högra axel och dricker en öl
En ung flicka blandar något gult i en skål.
En kvinna med brunt hår har en silverring på fingret.
En tjej i röd skjorta sitter med en laptop i knät.
Ett litet barn klättrar upp för en grind till ett stängsel.
En cyklist jobbar på sin röda upp och ner cykel.
Två kvinnor är utanför och gör något med krukor, kastruller och skålar.
Kvinnan justerar ett barns ansikte medan ett annat barn står bredvid hennes leende.
Det här är en man, som har ett rep i är mun, och en baby ko upp i luften
En grupp katter sitter i gräset.
En dam på en gård håller en hund medan en annan hund hoppar
Spelare gör sig redo för ett laserspel.
En kvinna som bär shorts matar två lamor eller alpackor på ett fält.
Vit fluffig hund som springer i smutsen.
En man med blå hatt och blå uniform som jobbar på lite utrustning.
En kvinna håller upp en bit spets som bakom sina män i ponchos spela musik.
Två män talar också en kvinna utanför, det finns träd runt omkring dem och en byggnad i bakgrunden.
En ung pojke i uniform nummer 24 skriker under en fotbollsmatch.
En man, klädd som polis, med en mikrofon i handen och ögonen stängda.
Dennis Hopper verkar prata med Cristy Ally.
En man med glasögon som tittar ner på något i sina händer.
Barn leker och gömmer sig under höet.
Någon håller upp en orm med huvudet och svansen mot kameran.
En arbetare står vid vagnen och tittar på något.
Unga män är närvarande vid en religiös ceremoni i en tjusig byggnad.
En kvinna balanserar ett litet barn på höften.
En amish dam förbereder en Clydesdale-häst för en vagn.
En man håller en kalv medan han slickas av en annan ko.
En man vinkar mot kameran och håller i en pinne med en trähög.
Två man spelar ett spel och stör.
Två fotbollslag spelar och en håller bollen igång medan det andra laget springer efter honom.
I ett vetenskapsmuseum som tittar genom ett teleskop.
Två motståndare fotbollsspelare med en i svart ta itu med den ena i vitt.
Ett litet barn som hjälper till att blanda något med en manuell mixer.
Två flickor och en förälder får ett studentrum i ordning för skolåret.
Två män som arbetar med jordbruksutrustning som dras av två hästar.
En ung svart flicka kommer ut ur badrummet inlindad i badrock och handduk.
Flera tonåringar röker och dricker på natten.
En ung flicka med overaller och galet hår sitter på ett grönt fält medan du äter ett rött och vitt objekt
Flera personer inspekterar de varor som visas i detta tält.
Man med svart hatt, vit skjorta och sandaler, lägger tegel på en byggarbetsplats.
En mycket leende baby som sitter ner i en randig jacka på en säng.
En dam klädd i rött skrattande med en dam klädd i gröna hålla tallrikar mat i sina händer.
En pojke och flicka är på en blå studsmatta.
Folk sitter runt ett bord med en röd duk som har mat på sig.
En man med slips pratar med två kvinnor.
En kvinna med grått hår tar en bild medan en man står bredvid henne.
En man visar en yngre flicka hur man dyker medan man tar itu med vågorna.
En kvinna med glasögon, bär blå jeans håller ett spädbarn medan pekar upp.
En kvinna knäböjer nära lyktorna medan en liten pojke leker i sanden.
En man som håller ut en deflaterad fotboll till en grå hund.
Två flickor klädda i vitt och en klädda i brunt.
En man i kostymjacka med ett gratis ordtecken.
Man tittar genom ett teleskop i en stad.
En man och ett barn under vattnet i en simbassäng som håller andan.
En liten flicka som planterar sin första blomma i sanden.
En ung pojke klädd i vitt och en skjorta läser "85" är i luften, gör en kampsport sparka.
En sångare i rampljuset poserar i sin läderjacka.
En mörkhårig kvinna som är dragen i en grå duk tittar ut ur en trädörr.
En pilot kör ett litet motorflygplan.
Barnet i randig skjorta balanserar mellan träräckena.
Tre arbetare målar utsidan av ett hus på byggnadsställningar.
Denna bild har en kontrollbord med fyra dryckesglas och ett askfat.
Färgglada Bollywood dansare i aktion på en scen.
En man, som bär en skjorta och en lungi, bär halmstrån på huvudet över en åkermark.
En man i blå skjorta står på stranden och kastar en sten.
En man med en floppig kockhatt håller i en kryddflaska medan han tittar över axeln som om han pratade med mannen bakom sig.
En vacker uppsättning färger visas från en dansare.
En stor fontän med flera personer som sitter på höger sida.
En man sjunger in i en mikrofon.
Den lilla flickan i poolen bär en röd baddräkt.
En visselpipa med vissling i munnen bär en bricka full av mat upp för trapporna.
En svart man i randig skjorta står och äter ur en kopp och håller i en gul vattenflaska.
Hunden springer genom skogen.
En man i den amerikanska flaggan simmar under andra vid en bassäng.
En kvinna i rött står med andra människor utanför.
En skjortlös sångare på en konsert framför en jublande publik med armarna uppe i luften.
En man tittar på sin kamera
En ung flicka slår en Scooby Doo pinata medan andra ungdomar och en vuxen observerar.
En kvinna i röd prickig klänning sjunger in i en mikrofon.
En man på en cykel och i bakgrunden en man utför ett trick på en skateboard.
Två barn ritar på väggen med kritor.
En grupp män och kvinnor som har ett möte utanför ett lager.
En gul hund fångar en frisbee i luften.
En man står på toppen av en stor höhög som dras i en vagn av två hästar.
En ung pojke som rider i en gunga.
Detta verkar vara en arbetsplats eller forskningsplats, möjligen en gård, men en mycket fuktig en som har några funky ser grön mögel krypande upp för väggarna.
Ett barn sitter ute i gräset.
En kvinna med blommor pratar i telefon bredvid en kvinna i bröllopsklänning.
Tjej med kort hår sjungande.
En vit man med blå skjorta står på scenen och sjunger en sång, hans svarta gitarrist står bakom honom och ger musiken.
En kvinna jagar två får med en kvast.
3 söta små flickor med något grönt i händerna.
En ung pojke i en hög med löv.
En liten pojke i svart t-shirt leker med en leksak NERF pistol.
En blond hund skakar vatten bredvid en sjö.
En leende man med en gul hård hatt kikar ut från ett manhål.
En man som pratar i en mikrofon med en kvinna som står bredvid honom.
En person på en balkong står bredvid några kläder som torkar på en linje.
Små flickor som har en födelsedagsfest som förklädes av en man.
En äldre man klädd i svart liggande på en grå möbel.
En kvinna med blå skjorta och örhängen.
En färgglad klädd man kör sin lika färggranna cykelrickshaw nerför gatan.
Ett barn som använder en dammsugare på köksgolvet.
En dansare i en levande rosa klänning som snurrar runt.
Detta foto är av olika individer som tittar genom teleskop i en plaza.
En pojke springer med en mycket liten fotboll på en asfalterad gångväg.
En Goalie i gult håller i en fotboll med en spelare i blått bakom sig.
En svart hund i vattnet med en tennisboll i munnen.
En ung flicka som gärna springer genom en park och håller i handväskan och leksaksbarnet.
Tre kvinnor i svarta rockar pratar och skrattar i ett konstgalleri.
En grupp vuxna sitter runt ett bord och spelar ett kortspel.
En dam skär en tårta medan den andra håller en tallrik med andra plattor staplade framför henne.
En man som bär en grön skjorta på banan driver upp en jetliner.
Lilla flicka i en blå och gul rutig outfit och blå hatt springer längs stigen.
En man gör sig av med vätska som finns inuti kartongbehållaren.
En person i en grön skjorta sitter på marken nära ett staket, med frukt utlagd nära henne.
En dykare står, böjd över på stranden.
En kvinna som sitter vid rosa blommor och hänger upp tvätten på en linje.
Den svarta hunden springer om vattnet med en rosa boll.
Tre barn och en man spelar volleyboll, barfota i sand.
En brun hund och svart hund födosöker i lite penselland.
Barn med lila skjorta och blå jeans är ovanpå en brun häst.
En kvinna med glasögon sitter i en stol och virkar.
En flicka som bär en pappershatt öppnar en present inslagen i rosa omslagspapper medan andra tittar på.
Två personer klättrar upp för en bärbar bergvägg
En kvinna i gult och blått hoppar baklänges över en bar.
En kvinna i en livsmedelsbutik läser över en lapp.
En publik tittar på när en stor man håller på att krossa något med en gummiklubba.
Grant var beredd att träffa sin golfboll medan hans caddy och målvakt väntade på honom.
En man i en lysrörsväst visar upp en modell av en byggnad vid ett möte.
En vildhund springer genom öknen.
Flickan sitter vid disken mellan hinken med blommor och pappkartongerna.
En man fiskar nära några vita vågor.
3 manliga cyklister stirrar på vänster sida av bilden.
En grupp på cyklister med sina cyklar på en parkeringsplats
En grupp manliga cyklister pratar utanför en bar med sin utrustning sittande på marken.
En flicka cyklar på en stig nära ett gäng träd och ett hus.
Två cykelcyklister rider sina vägcyklar genom en statlig park fylld med campare och andra cyklister.
Mannen i grå skjorta vilar en cykel mot ett träd.
Två män och en kvinna som står längst ner på en klippa.
Ett par klädda för en formell händelse poserar tillsammans.
En man i mustangskjorta gör sig redo att kasta en kniv på en tävling.
En hane och en hona vandrar i skogen.
En ung flicka bär kostym och lägger handen på hakan.
Cheerleaders kastar ut varandra i luften genom en fotbollsplan.
En ung flicka sitter på en blå bänk och dricker ur ett sugrör.
Två män i vita kostymer och glasögon med en drink.
En bicyklist i vita och svarta tights dricker framför en mini van.
En liten flicka i en rosa tröja använder ett teleskop på natten.
En äldre kvinna står vid skivspelare när en annan kvinna vänder på kameran.
En man i röda byxor som jobbar på sin cykel med en skiftnyckel.
Unga människor står i spray från en fontän under en molnig blå himmel.
En kvinna i orange utstyrsel böjer sig baklänges.
En kvinna som bär glasögon sitter vid ett bord och löder ett föremål.
En fiskare med en båt full av fisk.
En ung man som bär en rutig skjorta sjunger in i mikrofonen och spelar gitarr.
Män och två barn fångar fisk med nät.
En man i grön skjorta och blå jeans säsonger kött som det lagar kött på en grill på en bakgård.
Två hantlangare målar om eller rengör en tegelvägg.
En konstnär, bär blomtryck shorts och vit t-shirt, avslutar ett projekt med ett asiatiskt tema.
En man på en cykel körde just på en jordramp och är mitt uppe i luften.
Två pojkar leker med en leksaksbil.
Barn i ett klassrum som lär sig och är kreativa.
Män i vita och låga dräkter går med en stor fackla.
Deltagarna, klädda i långa vita tunika, på Burning Man Event poserar för gruppbild på kvällen.
Eleverna sitter uppradade på trappan medan de väntar och kollar sina elektroniska enheter.
En grupp människor deltar i en ceremoni.
Några ungdomar spelar ett kortspel
En grupp tonåringar plockar växter i en trädgård.
En pojke i rutig skjorta drar en vagn full av växter.
I detta foto finns det tre tonåringar som spelar fotboll.
En cykelförare glider nerför kullen mot en flagga, medan åskådare tittar längs den trädkantade vägen.
En fotograf skjuter en snowboardåkare i luften.
Detta är ett klassiskt café i europeisk stil, med en kvinna som står bakom disken och gör kaffe.
Klädd i sitt lag uniform av gult och svart han spelar fotboll.
Ett fotbollslag av unga pojkar som bär gula och svarta randiga skjortor är glada, när ett barn kramar en vuxen.
Barn som deltar i karateklassen.
Pojkarna är i karateklass idag.
Sex barn plaskar i en vattenpark utomhus.
En flicka med blå glasögon på huvudet gör ett ansikte medan hon ligger på gräset.
Singer fastnar i en hög ton och bryter en stämband.
En man i jeans overall och en röd skjorta gör jättebubblor för förbipasserande.
Sex musiker spelar sina olika instrument.
En barfota kvinna, nära en vattenförekomst, slår till mot en kampsport på hösten.
Poliser på hästar stannar av en grupp pojkar.
En kvinna som bär en tanktopp tänder en cigarett medan hon sitter med en annan kvinna.
En ung pojke hoppar fötterna först in i en inomhuspool.
En liten flicka klädd i mörka färger står på en klippa med utsikt över en stor damm vid parken.
En man och en kvinna i en stor röd klänning som dansar.
En man i mörk utstyrsel svingar en tennisracket, medan tre män i bakgrunden tittar på.
Några män sitter på soffor och spelar brädspel.
En man med blå mössa med vit långärmad skjorta och blå byxor spelar golf.
Tre män är på väg ut ur höet.
Ett fordon kommer över toppen av en kulle.
En kvinna drar en vagn med två pumpor i.
En grupp på sex personer sitter i ett möte och samtalar med varandra.
En man som håller två påsar i is kommer in i ett hus.
En far som spelar en sång på sin gitarr för sin son.
En pojke hukar sig bakom några små stockar och spelar paintball.
En man med läskig ansiktsfärg som bär en kroppsdräkt är fri att falla.
Flicka poserar på kanten av en veranda.
En tonåring sitter bakom en kartong och ler mot kameran.
En ung flicka slickar en tallrik och har tårta över hela ansiktet.
Den vita båten på vattnet har stannat.
Folk som jobbar på blommor i ett blomsterstånd.
Fyra män som bär t-shirts och spelar musikinstrument uppträder i ett band.
Barn leker badminton på gräsmattan.
En person sitter på en stor klippa medan en annan står i närheten
Lilla flicka kramar och bedårande katt
En man i orange skjorta använder en Mac-dator.
En man som talar in i en mikrofon med fingrarna i en nalle björn nos.
En man med väst och tan khakis shorts står ovanpå en bil.
En man sitter vid en bank av datorer medan han bär ett headset.
En man med mustasch och svart skjorta spelar saxofon.
En kraftigt påhittad brunettkvinna sjunger in i en mikrofon.
En kvinna i jeans och en grön t-shirt hoppar framför en silverstaty utomhus.
Två svarta hundar leker tillsammans på en gräsmatta
Två uppsättningar gatuartister uppträder för en grupp på tre på gatan hörnet.
Tre personer står vid några träd.
En sittande publik tittar på en man, bär en röd skjorta och svarta byxor och hängslen, lyfter en annan man, bär en mask, i luften.
Fyra barn som leker på en tältliknande struktur
Arbetare som gör sig redo att börja ett kvällsskift i ett närliggande företags komplex i staden
Två flickor håller i vattenkoppar medan de går bredvid ett taggtrådsstängsel.
En Pee Wee liga fotbollsspelare bär en lila jersey navigerar fotboll förbi motsatta spelare i vita tröjor.
Folk sätter upp stolar utanför på en parkeringsplats.
Fyra personer bär vitt är på en liten båt med andra båtar och nedslitna hus bakom dem.
En äventyrlig man navigerar genom djungeln med en lång käpp.
En collie leker med en vit boll i ett fält av grönt gräs.
Fyra män i mörka skjortor är på sina bärbara datorer.
Människor använder längst till vänster av tre rulltrappor, som är inneslutna i en avlång tunnel.
En man som spelar saxofon på gatan kanske vill ha pengar.
En man i svart skjorta håller i att spela musik på en gata.
Mannen i den vita hatten sitter vid bilderna.
Mörkhårig vit kvinna, bär en vit t-shirt och jogging byxor rakes blad
En liten blond tjej i gult skratt och springande.
En man med mohawk, skägg och skinnjacka sitter med en flicka med rosa mohawk och glasögon.
Folk går nerför trottoaren.
En man med en axellängd fram på scenen och håller en mikrofon med "Pop! Tech" skylt i bakgrunden.
En äldre kvinna jagar sitt barnbarn på en restaurang.
En person sover under ett bord täckt av en gul filt.
Det är många killar som springer tillsammans utanför.
Ett litet barn i en prickig tröja hänger upp och ner på en trädsving.
Barn ser på när en man dansar.
En hög vinkel vy av tre manliga musiker som uppträder i en mörk miljö med gitarrer fastspända på dem och en xylofon.
Fyra personer står nära skyltar och läser dem.
Många människor utforskar en konstinstallation på ett torg i staden.
En upplyst flicka stänker runt i naturligt vatten.
En kvinna med en svart jacka som sitter ner medan hon spelar piano.
En man som tittar genom ett teleskop med sin son.
En liten pojke är våt från att leka och skrika från strömmande vatten medan hålla en leksak valp.
En grupp människor i en stam går tillsammans.
En man gör en volt i luften från en sanddyn.
Arabisk kvinna köper frukt på marknaden.
En äldre man som skär en tårta för två flickor som sitter vid ett bord.
Två flickor med hästsvans rider på en nöjespark.
Ett litet barn använder en mixer på några ägg med någon annans hjälp.
En grupp människor som försöker plantera ett nytt träd.
En fotograf knäpper ett snabbt foto av en gul sportbil.
En flicka gör en kullerbytta mitt på ett gräsfält.
En kvinna med långt hår, glasögon och långärmad skjorta sitter vid ett bord och ler.
Två kvinnor och en ung man spelar ett spel runt ett bord.
En man och hustru utforskar en grön skog.
En blond-hårig kvinna med glasögon knäböjer bredvid en svamp i ett kraftigt vegeterat område.
Damen i rött sitter framför fontänen.
En musiker spelar en xylofon för en massa barn.
Två kvinnor som bär matchande huvudbonader säljer sitt goda på en marknadsplats på gatan.
Två män använder ett solteleskop för att titta på solen.
Ett gäng människor minglar på en mässa där det finns bås med flaggor av länder draperade över väggarna.
En pojke rider sin skateboard i parken.
Två kvinnor sitter vid ett bord, den ena tittar ner och den andra på en bärbar dator, med en banderoll som säger sweden i spanska bakom dem.
Två män vid ett bord diskuterar pappersarbete.
Två män i ett klassrum framför en vit skärm.
En man pratar och håller i ett papper.
En person åker skidor nerför en brant snöig kulle.
Två män med våtdräkter som rider på surfingbrädor.
En ung man i blå skjorta med vita shorts volleys en tennisboll.
En hund hämtar en tennisboll ur en vattenpöl.
En svart valp leker med en apelsin på ett heltäckningsmattat golv.
En hund som hoppar över ett stängsel.
En vit hund med mynningar på gräs framför träd.
En kvinna som läser en bok med matte.
Fyra män, klädda i vita overalldräkter som förhindrar infektion, är i ett rum med mekanisk utrustning och en stege.
En grupp vänner eller familj hoppar samtidigt för ett porträtt på semester.
De mörkhåriga barnen ler mot kameran medan en av dem sticker ut tungan.
En pojke med blå ansiktsfärg suger i tummen.
Kvinna klädd i vitt, sitter framför en stenvägg, spelar ett stränginstrument.
En man tittar in i ett teleskop.
Barn vänder sig till en folkmassa på rött tegel.
Unga svarta barn som dansar med tre som gör en pyramid.
En grupp på fyra flickor träffar en grupp äldre kvinnor.
En man i en orange mössa som står ovanpå en spetsig sten.
En brun hund med sele jagar en röd boll.
Två män som häller smuts på ett fält.
När en man går nerför gatan sveper en duva bakom honom.
Två män brottas vid en match medan åskådare tittar uppmärksamt.
En ung man utför ett rullskridskohopp framför en glasbyggnad.
En skidåkare hoppar över en lucka.
En clown i röda rutiga byxor och en rosa hatt sitter framför ett tält.
En svart hund bär en hink i munnen.
Cyklisten ler mot den våta hunden som slappnar av framför huset.
En ung kvinna skålar i UV-miljö.
En man knuffar två barn i en stor vagn medan en liten flicka springer bredvid dem.
Två barn arbetar med ett projekt med kvinna.
En man som bär glasögon och en trasig kostym spelar en Jaguar elgitarr och sjunger med ackompanjemang av en trummis.
En man i röd rock och svart hatt spelar trombon.
En asiatisk familj på fyra sitter runt ett kort bord.
En liten flicka med långt hår som flyter i en färgglad forrest.
En man som fiskar från en strandpromenad kastar sin fiskespö över räcket.
Ett ungt köp rider sin skateboard utanför på en ledstång.
En flicka står på en fot med en hand i luften.
En man i Elmo t-shirt cyklar genom skogen.
En hund i koppel sätter framtassarna på en bar.
En grupp människor, mestadels i orange och svart, går omkring under gnistrande.
En kvinna i svart klänning ler framför en silverbil.
Mannen med grön tröja och jeans faller från en stege när tre män tittar på.
Barnen framför byggnaden leker med en bubbla.
Vissa väntar på en busshållplats
Folk svingar på en röd, metall nöjespark rida framför några träd.
En kvinna i blå skjorta tittar in i ett skyltfönster.
En liten flicka i hatt och röda byxor balanserar på linor.
En man håller en gitarr på scenen under en konsert.
En far och tre pojkar går ner i vattnet på stranden.
En sångerska som sjunger i en rökig bar.
Ambulansen passerar en man som bär bandanna och flicka.
En man i svart utstyrsel kastar upp leksaksbollar.
En grupp människor som håller i väskor står i kö för ett tåg.
Helikopter landar i fält med sjö i bakgrunden.
En leende kille med glasögon håller upp en annan kille med en blå skjorta och svarta byxor utanför.
En man är på en skateboard på en röd ramp.
Ett afrikanskt barn har en fot på pedalen på sin cykel och stannar för att titta åt vänster.
Det finns ett par människor sätta dekorationer på en häst och en person tröstar den.
Den unge pojken med fina byxor, ett bälte och en slips hoppar från trappan
Grundskola barn passerar basket i lag basketspel.
En kvinna ligger på en randig soffa på en gräsbevuxen gård i ett bostadsområde.
Två personer i en föreläsningssal håller i en plastfolie.
Det finns en affär i ett främmande land med en man bakom disken.
Gentleman i en rosa skjorta slår trummor medan en publik tittar på.
En man med ett dystert ansikte tvingar sig själv att äta en ovanlig mat med ätpinnar.
En man och kvinnor steppdansar för en publik.
En liten pojke i en röd jacka står mitt i skogen.
Ett band som uppträder i hörnet av gatan.
Skateboarder gör en kick av en upphöjd plattform på en trottoar.
En man paddlar en kanot tillsammans med en hund.
Man med lila hår och en blå skjorta som fixerar ett vakuum med en annan vit man, som är äldre.
En man kör sitt bagage förbi ett fönster fullt av blommande blommor.
En dam som står på ett utställningsbord för en ringkastning.
En flicka i rosa och man i svart paddla genom vatten.
Ett par unga män sitter på en stoop i ett nedslitet område; en verkar vara metallbearbetning.
En man uppträder för en grupp framför ett vitt hus.
Män som går på stadens gata med en gul buss och två FedEx fordon i bakgrunden.
En man och en ung flicka som simmar.
En grupp barn tittar på en skulptur i ett museum.
Tre män spelar långa trummor på en scen.
En hund har en orange boll i munnen.
En kille som rider motocross i smutsen.
En grupp människor går uppför en ramp en molnig dag.
Afrikanska män dansar medan de bär en blandning av traditionella och västerländska kläder.
En äldre man i svart skjorta sitter med tre små barn utanför.
Man med stormtrupper huvudbonader på affärer för godis.
Tre afrikanska kvinnor dansar i infödda afrikanska kläder medan en grupp människor tittar på.
Man sover på en gammal soffa i en gränd.
En man som går mot en vit glassbil parkerad på gatan på natten.
En flicka tittar på en insekt på fingret och ser rädd ut.
Ett ställe som ser ut som en fallskärmsanläggning folk sätter på hjälmar.
En man med en fiskespö som står på en strand.
En tatuerad kvinna spelar gitarr och sjunger medan hennes band står där bak.
Två flickor i kjolar som ler i en park.
Två kvinnor i rosa overaller poserar bredvid ett vitt fordon.
Asiatiska män och kvinnor som sitter på blå plastpallar äter.
Ett tremannaband spelar på scenen.
En hund som springer genom vatten.
Denna hona med tatueringar sticker ut sin genomborrade tunga, medan hon håller i en ölburk.
Kvinnor sminkar sig medan de pratar och pratar i telefon.
Ett barn rider en enhjuling längs en stig intill en kvinna som går en hund.
En svart hund leker runt nära ett vattenfall.
En man står framför en torktumlare i en tvättomat med båda händerna i en soptunna eller korg.
En man som bär svart hatt är ovanpå en travhäst.
Springer snabbare än en fortkörningskula och är på väg att köra om den vita sedan.
En man i kostym rider en brun häst.
Ett lugnt gathörn med en man som sitter på en pall och tittar på något på en liten plattform.
Killen i en blå skjorta vänder hamburgare och korv på en utomhusgrill.
En man som bär glasögon med hjälp av en spatel för att lyfta en hamburgare från grillen.
Två personer som gör sig redo att servera mat till andra.
Två män arbetar med keramik i ett rum med keramik på alla väggar.
Flera män drar ett fiskenät upp till stranden.
En man i militärdräkt pratar på en bärbar telefon.
Hund sitter på ägare knä sitter framför datorn
En asiatisk man som försöker reparera en grön cykel utomhus medan två andra asiatiska män väntar.
Familjen dansar på sidan av en sjö vid solnedgången.
En flicka i svart kjol och blå klänning vattnar blommor.
Många barn samlas runt ett bord fyllt med mat.
En flicka i en långärmad t-shirt med flerfärgade ränder, och svarta byxor, äter en topping från en hemmagjord pizza hon förbereder.
En ung blond pojke äter tårta med en sked.
En unge med en blå Mohawk spelar fiol
Barnet är fascinerat och fascinerat av hans bild i vattnet.
En liten pojke som bär badbyxor leker i havet.
Två barn glider nerför en vattenrutschbana på en uppblåsbar flotte.
Två indianer säljer chips till fotgängare som gatuförsäljare.
Hemlös man som ber om pengar med hjälp av humoristiska tecken.
En äldre man i rock och stövlar förbereder en nyfångad fisk.
En man på en mikrofon som spelar piano och tangentbord.
Ett barn gör ett handstånd vid kanten av en strand.
En grupp män på en båt som är tipsad med hjälmar.
En ung pojke i en tom hall med två andra i bakgrunden.
En äldre herre som visar stolthet när han visar upp sin trädgårdsskörd.
En svart man som håller i ett hök.
En man på en stege som gör något med torkade växter.
Två män, en i svart skjorta, den andra i jacka, staplade vete.
En kvinna i en trenchcoat som anropar en taxi för en åktur.
En brunhårig pojke i badbyxor vänder sig baklänges över en simbassäng.
Ett litet barn plaskar i en grön och gul vadderingsbassäng
En man som bär solglasögon och bär röd väst står framför en röd helikopter.
En flicka i rosa klänning leker med en hulahoop.
En kajakpaddlare i vitvatten forsar mellan två stenar, och en åskådare på en stenig strand tittar.
Två barn forsränning på en sjö.
En liten flicka sitter i ett metallbad fyllt med vatten.
En man på en moped kör genom gatorna i sin stad.
En person som bär en mikrofon har ett rött täcke över huvudet när han går framför ett svart täckt bord.
En Cirque de Solei-artist visar upp sin imponerande styrka och balans.
En flicka dras av ett snöre medan hon sitter på en flotte.
Två pojkar leker med en skadad fotboll.
En pojke i en bilstol sover och gråter.
En ung flicka i glasögon och träningsoverall svänger ett racket.
Ungdomar med matchande frisyrer poserar för kameran under ett vitt paraply.
En liten flicka i gul skjorta med en stor snigel.
En ung blond hona tenderar till en liten valp utomhus.
En man i orange skjorta som klättrar på stenar.
En man med glasögon och en grön skjorta blir kysst på kinden av en biffig get.
Många människor sitter nära Space Needle.
En person på skidor rensar ett hopp i ett vackert berg täckt av snö.
En liten flicka är utanför och håller i en snöboll.
Ett band sätter upp en ljus show och en föreställning framför en publik.
Fotbollsspelare tar betalt mot varandra på det gröna fältet.
En kvinna som cyklar förbi en bil och en grupp människor på en trottoar.
En liten pojke som knuffar sin trehjuling mot bollar som ligger i gräset.
Mörkhårig konststudent som arbetar med ett projekt medan han ställer sig upp.
Tre arbetare lyfter en röd säck medan en annan sitter på en flytande docka.
En man ler för att ta fotot medan han arbetar.
En ung svart flicka ritar färgglada blad på papper.
En ung man som tittar på himlen genom ett personligt teleskop på kvällen.
En man använder sin dator när han sitter vid ett skrivbord.
En motocross ryttare, rider längs en grusväg på en solig dag.
Mannen sveper med en röd kvast.
Två barn, en pojke och en flicka, i luften ovanför en studsmatta.
Ett stort plan som håller på att monteras ihop.
En dam målar många lådor.
En stor grupp människor höjer sina händer vid ett möte.
En ung pojke leker med leksaker bredvid en kvinna som ligger på golvet.
Den lille pojken njuter av föräldrarnas sällskap.
Människan sopar skräp från vägen med en bunt kvistar.
En skateboardare bär blå jean och en grå skjorta utför ett stunt längs en graffitifärgad vägg.
En man väntar vid en busshållplats bredvid en lastbil täckt av graffiti.
En man flyger genom luften över en stor kanjon.
En man som flyter omkring på vattnet och tittar på något vitt i sina händer.
Barnen åker båt i vattnet.
En man med en orientalisk hatt som plöjer ett fält i en blå skjorta.
Två flickor i kostym sitter på en trottoar.
En gammal kvinna i ett solbelyst rum slingrar grova garn till bollar, de färdiga garnbollarna placeras i en hög till höger om henne.
En grupp människor köper mat från en säljare.
De tre rockstjärnorna är medlemmar i ett band som spelar på en konsert där färgerna rött och svart är framträdande.
En fotbollsspelare springer mot en annan spelare.
En kvinna klädd i en svart jacka som vilar på en hylla på dryckesavdelningen i en affär.
En man håller i en pinne medan tre hundar tittar och hoppar.
Tre kvinnor arbetar på ett fält, medan fyra barn och en dam håller en barnklocka.
En kvinna i en flerfärgad skjorta gör en hängmatta.
En man bär en tröja och jeans denim spelar gitarr medan en kvinna spelar trummor
En nunna tar en bild utanför.
En man i blå skjorta går en cykel laddad med en stor låda på baksidan.
En pilot städar ett fönster på flygplanet.
Fyra män står nära ett brödstånd utanför medan en av dem tar en tugga.
En leende kvinna bär två korgar fulla av råvaror på en bambupåle.
En grupp musikaliska artister spelar och en skara människor finns runt omkring dem.
Två män som tillverkar kläder i ett tredje land.
Köpmannen gör i ordning sin monter med välsmakande etnisk mat som skall säljas på marknaden för utomhusbruk den dagen.
En pojke klättrar på en hög av trä trots en skylt som förbjuder det.
En person, klädd i hatt och lila tröja, målar en hamnscen.
Två barn är klädda som pirater.
En person duschar i ett mörkt rum.
Två barn i piratdräkter slåss med sina svärd.
En pastor och en ung flicka framför katedralen.
En man arbetar på ett ofärdigt tak.
Flera personer håller moppar stående runt två gula mopp hinkar.
En plysch tecknad maskot poserar med en ung flicka.
En ung skidåkare njuter av backarna med stolliften i bakgrunden.
En snowboardåkare som gör ett stort hopp gör ett trick på ett högt berg.
Det finns tre kineser som är på en paus från fisket.
De två flickorna njuter av att åka pulka i snön.
En brun hund och en svart hund på en grusväg.
Folk går genom en gata på natten.
Två asiatiska män som arbetar på sidan av en gata med parkerade bilar.
Unga par gifter sig i en park omgiven av träd.
En asiatisk man cyklar nerför gatan, där blommor och andra fordon finns.
En flicka som leker är en hög med färgglada bollar.
En pojke i en blå skjorta tittar på en kvinna som bär en mångfärgad klänning medan ett annat barn ser åt motsatt håll.
En man bär kostym och kör en vagn.
Hunden sover ovanpå sängen täckt av det blå lakanet.
En båt som heter "ELOIN" flyter på vattnet.
Ett blond-hövdat kvinnligt barn som leker med leksaker på en lila yta.
Två flickor utövar yoga i en park.
En ung pojke i en blå skjorta som iakttar en skör boll som hänger från ett rep.
En gammal man och en ung kvinna dansar tillsammans medan åskådare ser på.
Pojke på skateboard ridning framför höga betongstaty med brons staty på toppen.
En man sitter med fiskestolpar nära en vattensamling.
Sju personer, mestadels i vita skjortor, dansar i ett rum med en röd vägg.
En man har en skylt som erbjuder sig att byta en dikt mot en fotbollsbiljett.
En mörkhårig gentleman med mustasch och tröja trycker samtidigt på knappar på en gammaldags datormonitor och tangentbordet.
En bebis tuggar på en leksakslastbil.
En man som spelar elgitarr framför en bakgrund med flygplan.
En kvinna i gul blus som rakar huvudet på en annan.
En man som deprimerande glänser ner när han ser en majoritet av sitt hår falla ner på golvet vid frisörerna.
Fyra personer bär snöskor hoppar på ett snöigt berg med träd i bakgrunden.
En basketspelare tar ett fult skott som sina lagkamrater och motståndarlaget klocka.
En man med en stor kraftborr står bredvid sin dotter med en dammsugare slang.
Ledarsångare för ett band håller i en mikrofon.
En man bär en svart hjälm och är på en svart skateboard.
En grizzly-liknande man med stort skägg spelar tangentbordet med en kvinnlig bandkamrat som spelar gitarr.
En gammal gitarrist utan skjorta pekar, svettas.
En man i blå skjorta och en man hjälper cyklisten medan mannen i grå jacka klockor.
Man försöker plocka upp motvillig flicka på gatan.
En tjej som bär baddräktströja bär ett tecken för att ge gratis kramar.
Den stora dansaren slungar runt håret.
En pojke i badbyxor plaskar i en simbassäng.
Två män och en kvinna som sjunger och spelar instrument på en scen.
En pojke hoppar ner i vattnet med en boll i handen.
Män klädda i arbetsutrustning bedömer ett dräneringsområde.
En blond tjej poserar för en bild på Kerry Park i Seattle.
Tre män nära vattnet med gula västar och hjälmar.
En kille med en orange, grå och blåjacka som drar en kärra nerför en trottoar framför en väggmålning på en byggnad.
En man i randig topp skriver på en svart tavla.
En äldre man som joggar på ett löpband gjort av Life Fitness.
Detta kan vara en jobbmart eller möjligen en röstningsstation.
En svart hund närmar sig en gyllene hund på stenig strand.
En kvinna i blå snödräkt åker skidor, medan hon släpar ett träd bakom sig.
En kvinna på skidor som går uppför en kulle och bär en tall.
Lastbilschauffören stannar för en fotomöjlighet.
En liten flicka i rosa pyjamas leker med en leksak hus som hennes mormor vakar över henne.
En kvinna i en tryckt utstyrsel bär en bricka på huvudet.
En person i smutsiga kläder skär sten och skriver något i Urdu
Ett antal personer på en pir är silhuetterade mot solnedgången.
Folk utforskar en stad med sina kartor och kameror.
Tre street hockeyspelare spelar ett spel.
En man som håller i en resväska går ensam mot en rulltrappa i ett svagt upplyst område.
En hund hoppar över baren.
Människor som håller parasoller över huvudet går upp för en trappa bredvid en rulltrappa.
En kvinna sjunger och spelar gitarr.
Två personer sitter på en bänk med sin hund bredvid en vattensamling.
Två barn som ligger på marken ler mot varandra.
En pojke med röd hatt chockad av att en lekplatsleksak snurrade.
En man som tar bågar på vägen.
En ung afrikansk man som håller en penna i varje hand och studerar en bok medan han sitter nära ett öppet fönster.
Kvinnorna i de blommade byxorna gör trädgårdsskötsel.
En man böjd över i en skog bär en röd skjorta och blå jeans, knackar träden för lönnsirap.
Många människor flyger färgglada drakar på stranden.
Kvinnan i den blå rocken pratar på mobilen medan hon hänger upp bensinpumpen.
Jermaine från Concords flykt lär ut matte i ett främmande land.
En målare sitter på en gunga för att hjälpa honom att måla väggarna i en byggnad.
En rullande nål tillplattande gulaktig deg.
En mager kille äter en smörgås medan han använder datorn.
Kvinnan sveper gatan med en röd jacka.
Ett gäng ungdomar som dricker på en bar.
Medlemmarna i Frälsningsarmén står tillsammans när man innehar ett instrument.
Två händer måla en bild med endast färg, cirkulära lock och fingertoppar.
Två unga pojkar brottas i en sandlåda.
En man i väst och slips spelar gitarr på trottoaren.
En lättklädd man spelar gitarr.
Gruppen arbetar med mikroskop och bär rena vita skrubber, hårnät och ansiktsmasker.
Tre personer sitter på en soffa inne i ett hus klädd varmt och den äldsta täcker de två yngre barnens ögon.
En man med solbränd hatt och jacka fiskar i gröna vatten.
Tjej på rosa skateboard bär svart jacka
En cellospelare och en violinist som gör sig redo för sin föreställning i ett elegant rum.
En närbild av en vit hund som dricker ur en pipa.
En kvinnas fiskespö är nedböjt när hon står på en båt i havet.
En hane i svart kostym och hatt som håller garn.
En arbetare använder en jackhammer på stenblock från en klippa, en soptipp står parkerad i närheten.
En byggnadsarbetare gräver ett hål på gatan medan en annan man tittar.
En grupp människor rider nerför en berg-och dalbana som verkar kallas "Cyclone".
Medlemmar i en bygggrupp diskuterar ett problem med ledningen.
Två byggnadsarbetare i orange västar rider i en bit utrustning.
Manlig vuxen utövar skateboard tricks på en skatepark.
En man i en gränd gör sig redo att kasta ett föremål upp till någon ovan.
En grupp människor trummar medan de sitter i en cirkel på ett gym.
En skadad fotbollsspelare på kryckor, bär en röd vit och blå uniform, ser mot himlen.
Folk går förbi gamla vita väggar med grå rutor.
Två kvinnor arkiverar i wrappers medan en man med en blå t-shirt ser på.
En hund som springer genom gräset.
Två killar i ett främmande land som lagar mat över en grill med folk som går runt dem.
En ung man tittar på foton på sin dator, sitter vid ett skrivbord.
En liten flicka lutar sig över ett litet stängsel och tittar noga på en ko.
En man lutar sig tillbaka i en stol och dricker läsk och äter.
Två män, en John McCain, och en kvinna som sitter i röda rullstolar bredvid en vit skylt med en blå bokstav D och en nummer 5 på den.
En ensam bodyboarder med en äldre man i bakgrunden
En man med glasögon i brun skjorta pratar medan en man med glasögon i grå skjorta lyssnar.
Man i shorts och t-shirt på väg att börja använda gliding träningsutrustning.
Två män på en pratshow tillsammans sitter i röda stolar.
En man målar en livfullt färgad stadsscen.
En grupp människor står på en gata med höga byggnader till varje sida av dem.
Folk går på en vacker dag i San Francisco.
En liten flicka gör ett fånigt ansikte medan hon håller en trofé utanför.
En klättrare i en gul hårdhatt ses mitt i klibben uppifrån.
Tjej med långt svart hår och vit hjälm, häller vatten från svart vattenkokare i muggar.
En shoppingplats med många människor.
Två ungar skyfflar snö och en sitter bredvid snöhögen.
Händerna med målade naglar avskruvande nagellack.
En man i blå dräkt lagar mat medan han är omgiven av tallrikar med grönsaker.
En bowlare ska kasta en grön bowlingboll nerför gången.
Två personer sveper i en struktur som har kolumner med bilder på sig.
En vacker ballerina med julljus runt kroppen.
En ballerina i en grönaktig och blå outfit hoppar under sin föreställning.
En kvinna och en man som spelar bowlingspel
En svart hund på en brygga som ska dyka ner i vattnet efter en boll
En svart hund på koppel som går i vatten
En kvinnlig vetenskapsman och en manlig vetenskapsman tittar på en bok tillsammans i ett labb fullt av växter.
En man i vit skjorta som sitter med en kvinna i en blå blus.
En ung man som använder en lövblåsare för att rensa höstsäsongen lämnar området.
En person som bär stora glasögon läser en orange inbunden bok.
Fem personer i blått räfsande gräs framför en vit byggnad med en blå balkong.
En grupp turister tar en tur på en häst dragen vagn.
Ett barn hoppar på en struktur täckt med mjukt material.
En gammal kvinna som bär solhatt och rosa blus undersöker ett gräsigt, träskigt fält.
Två små pojkar tävlar mot varandra medan en liten flicka tittar på dem.
En kvinna i solglasögon som fotograferar
En ung pojke sitter på golvet och försöker ta av sig stövlarna.
Kvinna med puffig jacka tittar på soppa objekt i en livsmedelsbutik.
En grupp unga vuxna män har monopol.
En kvinna bemannar en grill med lite kött
Folk grillar aktivt på grillar en solig dag medan andra står i närheten.
En man i blå skjorta leder barn.
En galen som sitter ner och borrar ett hål i en glasflaska.
En man med kort hår och ett barn sitter när barnet öppnar en present.
En man med skägg och väst dekorerar sin mantel med strumpor till jul.
En kille som fixar en datordel och tittar på den som tar hans bild.
Två personer går i motsatt riktning över en tegelväg.
En ung pojke som bär glasögon arbetar med ett enkelt vetenskapsprojekt.
En liten pojke leker med en gul spade framför en julgran.
Fyra personer i flytvästar flyter på en flotte.
Två kvinnor står utomhus en vinterdag på landsbygden.
En kvinna med disk i smutsen.
Tre kvinnor vilar vid ett bord med blå servetter och kannor med vatten.
Äldre gentleman med långt hår talar in i en mikrofon.
En mörkhårig person i en gul topp sitter på vad som verkar vara ett flygel.
En ung pojke i en brun jacka som spelar piano.
En man som bär en rutig kortärmad skjorta och ljusbruna byxor hoppar högt i luften framför dimman täckta berg.
Två bruna hästar drar en släde genom snön.
En blond bebis ser en mörkhårig bebis tugga på en blå leksak.
En kvinna spänner fast ett vresigt barn i en bilstol.
En mångfaldig grupp människor som sitter på trappan och halva väggen framför en skola.
Två män sparkar fotboll på en strand.
En medelålders asiatisk kvinna på ett evenemang som visar en röd korsett för en publik.
En byggnadsarbetare står på en träbjälke och tittar ner.
En glad grupp människor ler för en bild på en restaurang
En grupp människor dricker kaffe och får lite arbete gjort.
En man i svart topp hoppar på en solig dag.
Många män i lila spelar trumpeter.
En man i vit Coca-Cola-skjorta och newsboy-hatt lyssnar på ett bandspel.
Grupp sitter på en gräsbevuxen kulle vilar.
En barfota kvinna i svett hoppar upp i luften med andra på liknande sätt klädda människor bakom sig.
Ett leende litet barn bär en kostym.
En man står ovanpå en elefant i vattnet.
En ung pojke tittar på en uppvisning av gummiankor.
Ett par människor går på en stig med en stad i fjärran.
Den lilla pojken går nerför kullen medan en äldre kvinna tittar på
Solglasögon som bär ung vit pojke står på ett fält av vita blommor och håller en fotbollsboll.
En polis på en motorcykel som pratar med två män på en kullerstensgata.
En pojke, klädd i svart och blå snödräkt och snöskor, ligger ner i snön.
Två personer bakljus med ljus himmel.
Den här tjejen sjunger inför många människor som bär en fin, moderiktig klänning.
En man och tre pojkar sitter på parkbänken
En skuggig man som tittar på de avlägsna kullarna.
Två små barn leker med färgglada leksaksbilar på golvet.
En kvinna i lila kläder som går längs trottoaren och bär en vit väska.
En träningsklass med deltagare som cyklar stationärt.
En man i lila och vit skjorta hjälper en man i en hustrumisshandlare med sin träning.
En förälder rakar ansiktet medan ett barn bråkar med håret.
En man målar en scen av en sjö och båtfolk medan en annan man tittar.
Två hundar biter varandra i snön.
En äldre man sållar vatten genom fingrarna när ett litet barn tittar inifrån vattnet.
En reklamtavla annonserar en semester på en nedsliten gata.
En grupp ryttare färdas längs en grusväg.
Tre personer klättrar upp för ett berg på skidor.
Snowboarder bär en orange jacka och bär en himmelsblå väska snowboards mot en tidigare rest spår.
En man knuffar en ung flicka på en scooter.
Två män som städar fönstren i en hög byggnad
En ung man som snowboardar på natten är mitt uppe i luften och gör ett trick av ett hemgjort skidhopp.
En man i ett badrum ser ut i spegeln och tillämpar rakkräm.
En åkare som maler ner en räls framför en latinbutik medan tre åskådare tittar på.
Två unga damer i en bar som dricker vin till en skål.
Fyra balettdansare i svarta kostymer uppträder på en scen.
En man i orange jacka faller ner i en snöig bergssluttning.
Två tungt klädda människor förbereder sig för att göra te i snön vid en lägereld.
Tre personer går genom snön.
En liten pojke står i dörren till en skåpbil.
Ett vitt och rött skepp fyllt med människor sitter i vattnet medan en rad andra gör sig redo att gå ombord.
En svart hund kommer ut ur en röd tunnel.
En stark kvinna i blå skjorta lyfter vikter med en maskin.
En kvinna som hoppar i en öken som ett område.
En skara människor står utanför med rockar och paraplyer eftersom det regnar.
En skjortlös man med en hund bredvid honom som pratar med en skjortlös flicka som slumrar på en bänk.
En hand som petar ur en svart tröja är att blanda ett ägg till en mjölbrun med en gaffel.
Ett barn drar en leksak genom en fontän med andra barn och människor som tittar på.
Tre män står i en polisbåt med många stenar bakom sig.
En dam applicerar svart naglar på ett klädbord.
En ung man i röd rock ler.
En grupp män från Mellanöstern som säljer småsaker på gatan.
En kille med långt hår och vinglas står nära två andra män.
En liten pojke i blå randig skjorta kommer nerför stora rutschkanan.
En brun hund hoppar när han tittar på en fotboll.
Fyra äldre män spelar poker på en uteplats.
En man med mycket rörmokares crack väger en sten, av någon okänd anledning.
Ett barn i en färgglad hatt inspekterar sin snöängel
En äldre man som använder ett mikroskop för att få mer finess i träbearbetning.
En man sätter gräs på en bil dragen av en gräsklippare.
En liten pojke med blont hår tar ett bad i ett litet blått badkar.
Ett band spelar musik i en ljusfylld scen.
En man i brun jacka sitter och arbetar på en detaljerad målning.
Tre personer står vid disken i en affär.
Två unga flickor sitter på marken och gör något av halm medan en liten pojke sitter mellan dem.
Man hoppar på sidan av vägen bredvid en bil full av vänner.
En kille som ler med en pinne i en färgburk.
Fyra killar i vita kläder är i en studio.
Ett litet barn står utan tröja i en mörk skog och håller en liten fågel i sina händer.
Hunden står i sanden nära havet.
En pojke står framför en skrothög som innehåller metallskrot och en skadad bil.
Kvinnan pekar på ett konstverk med glas som täcker det.
En pojke i baskettröja och svarta sportshorts står på ett ben på en gata.
En grupp män spelar fotboll i öknen.
En ung kvinna i blått bär en låda i ett ofruktbart rum.
En mycket ung flicka sitter i en livsmedelsvagn i närheten av en livsmedelsbutik deli.
En ung flicka leker med en leksaksbläckfisk framför sin julgran.
Tre barn leker med en grupp ankor.
Tre personer leker i snön med en skog i bakgrunden.
En sångare uppträder med sina bandkamrater som spelar gitarr och keyboards.
En pojke med åra går ut från surfingen och upp på en strand.
En kvinna skjuter ett gratiskast på en basketmatch.
Två barn hoppar på en säng, den lilla flickan är i svarta byxor och är mitt i hennes hopp.
En kvinna poserar för bilder med en staty av ett troll.
Ett gäng hipsters i bowlinghallen verkar reagera på chockerande nyheter.
Två kvinnliga basketlag tittar på spänning när basketen närmar sig korgen.
Tre personer står framför en flod vid en stad medan man kastar något i den.
En grupp människor hänger upp och ner på en berg-och dalbana.
En grupp på fem personer rider i en kanot i en flod.
En grupp människor rider i en hästritad vagn.
En liten pojke i polotröja äter något.
En brun hund hoppar ner i en damm.
En kvinna och barn står bredvid en stor brandbil.
En välklädd man håller en saxofon och går framför ett piano.
En ung flicka som bär en blå skidmössa och röd och grå tvåtonig jacka står mellan två bitar is.
En ung flicka med ett målat ansikte springer på en bakgård.
På ett fantastiskt blått tropiskt hav sitter en man i sin båt och lagar sitt fiskenät.
Två personer gräver marken av ett gäng båtar.
Det ser ut som om flickan gick och handlade och fick något från AVEDA-butiken.
En man som går sin hund på en korsning.
Fem personer arbetar längs stranden i ett asiatiskt land.
En person som står framför ett flygbesättningsmonument.
Fyra till fem ballerinor gör en dansensemble på scenen för massorna.
Stor hund försöker bita liten hund
Människor står nära vattnet med en båt på väg mot dem
En oförskräckt koflicka rider en mustang på rodeon.
Två herrar tittar på sina grödor strax utanför ett skogsområde.
Två unga pojkar tittar på någon på en skateboard.
En kvinnlig talare på SVA-teatern håller tal.
En kvinna och en cocker spaniel leker i snön.
En pojke i en röd hjälm träffar en boll med ett slagträ.
Ett barn får lära sig av en vuxen att rida på ett får.
En campingplats har etablerats bland träden och buskarna.
En man med grå skjorta klipper gräsmattan medan hans son gör samma sak bara med en leksak gräsklippare.
En person med skidmask, handskar och solskydd ligger på snötäckt yta.
En ung flicka och pojke på en åktur på en nöjespark.
Person som går genom snö lövlösa träd i bakgrunden
En kvinna och en man är på en självkontrollstation.
Två små pojkar i en kanotpaddling nerför floden.
Två kvinnor rider hästrygg över en gräsbevuxen kulle.
En person cyklar nerför vägen, medan en annan sitter i en båt på vattnet.
Två hundar utanför slåss om en röd Frisbee.
En grupp unga vuxna samlas för att framföra sång komplett med trummor och en gitarr.
En ung boll somnar i en kundvagn.
En kvinna med öronmuffar har ett papper som säger "verklig förändring" på omslaget.
En peloton av cyklister som rider längs en väg av tätt packade hus.
En pojke och en flicka tittar på ett blått Nintendo DS-spel.
En kvinna draperad och udda klänning, läser för publiken.
Två personer fiskar på en brygga med en lång slingrande bro i bakgrunden.
En byggnadsarbetare passar ihop metallrör.
En person som bär snöskor står i snön nära en bäck.
En kille som kör sin fyrahjuliga smutscykel medan han tävlar.
En man spelar gitarr på en scen, ljuset lyser bakom honom.
Ett hockeyspel har det vita laget mot det svarta laget.
Lilla flicka i jeans och en rosa skjorta vadar längs stranden.
En grupp människor väntar i liknande klädsel.
En man som bär hatt och förkläde provsmakar en smak av sjudande soppa.
En man målar sidospåret, av tidigare beige byggnad, vit.
En liten svart hund jagar ett stort djur i ett inhägnat område.
En kvinna kämpar med att svinga en hoe medan hon skördar på ett fält.
En ung asiatisk flicka i en tub topp håller ut sin kamera för att få en bild med sin vän som gör fredstecken.
En rödhårig kvinna ser förbi kameramannen.
En tjej i röd tank och jeans sover på en brun soffa.
En flicka står bredvid en hund medan hon lutar sig mot ett staket och står på marken.
En kille i morgonrock som sitter på kanten av en bubbelpool och ler.
En mycket svag kvinna håller i en gryta och några grenar ovanför huvudet.
En fullstor häst och ryttare styr en pint storlek häst och ryttare genom stallet.
Ett barn tittar genom kikaren på en båt medan hennes yngre syster väntar bredvid henne.
En flicka som tittar över axeln ligger i en rabatt och längs en gata.
Två kvinnor med sitt hår täckta samtal i ett kök.
En kort tjej i vit kjol, svarta stövlar och en grågrön jacka som bär en röd väska på trottoaren.
Två människor klädda som djur nära en folkmassa.
En pojke i svart viftar med armarna medan andra står bakom honom på ett fält.
Två kvinnor med kjolar som går längs gatan tillsammans
En ung man utan skjorta, som står under lila ljus, pekar mot himlen med båda händerna samtidigt som han håller en mikrofon i en hand.
En man som går längs och torkar golvet på flygplatsen.
Den svarta hunden och den bruna hunden verkar vara brottning.
En ung flicka svävar i ett metallbad i en vattensamling, medan hon håller i en orm.
En svart hund springer nerför en blå och orange ramp.
Grupp av längdskidåkare vandrar upp för ett berg.
Två personer i skidor, bär blå jackor, med ryggsäckar står i snön på ett berg nära en markör.
En liten barn hängande upp på lekplatsen
En brun och vit Sheltie hoppar över en räls.
Ungt barn som leker med en fotbollsboll i ett gräsbevuxen område.
Här är soldater i transport i ett fordon till någon plats, de är omgivna av andra soldater och utrustning.
En pojke i grå träningsoverall packar upp ett DVD-spel.
Två barn är på en enorm uppblåsbar rutschbana.
En man i en morgonrock blåser bubblor i ett badkar.
En kvinna med glasögon sitter på en gunga, på en lekplats med många träd.
Tre personer som cyklar på trottoaren.
En flicka i en tröja är i ett tempel med en mängd olika växter.
En man talar in i en mikrofon på ett konstgalleri.
Två hanar rider på hästar som jagar en ko på en röd träarena.
Fyra män uppträder musikaliskt utanför en byggnad.
En skara människor tittar på ett musikband som är under ett tält.
Fem personer sitter tillsammans och spelar instrument.
En två asiatisk kvinna som målar ett trästycke.
Två killar med snöskor som tar sig genom skogen.
Två män både bär cowboyhattar och ponchos rider hästar jagar en ko.
Tre män på hästar jagar en tjur på en arena.
En ung tonårspojke som krigar med en grön snödräkt hoppar över en uppsättning kraftledningar medan två kvinnor tittar på.
En man i en brun rutig skjorta har händerna på en bils strålkastare.
En kille som hoppar från en brygga ner i en vattensamling.
En postarbetare håller i en handfull varor som skall levereras.
Fyra musiker spelar sina instrument på gatan medan en ung man på en cykel står och lyssnar.
Tre män med trummor och tatueringar står nära en kille som spelar säckpipa.
En skäggig man spelar trummor i skymningen, och en man som sitter bakom honom spelar en elektrisk gitarr.
En kvinna är upphöjd på en soptunna och fotograferar.
En man som bär snöskor går nerför en kulle bredvid små orange flaggor.
Människor i snöigt klimat förbereder sig för att äta mat på tallrikar.
En parad av män håller röda och gula flaggor när de vinkar stolt.
Grupp av människor som står och sitter i ett fält av gräs.
Flickor som bär en blå klänning med ett tunt, långt, blått tyg medan en flicka ler och pekar mot kameran.
En kvinna går på trottoaren bredvid graffiti taggade väggar.
Polisen och brandmännen diskuterar vad de ska göra med den välte SUV som ligger i snön.
En blond hästsvansad kvinna och en gråhårig man samtalar medan han sitter på en restaurang utomhus.
En man i blå jacka ler tillbaka mot kameran, placerad framför en sjö eller stor flod på en klar solig dag.
Män förbereder ett segelfartyg vid en docka.
En kvinna som bär skridskor, hjälm och kuddar, hoppar upp i luften.
En man i blå skjorta och byxor står framför en stor skylt som visar en jak.
Två personer i en båt, en en röd skjorta och en i en grön skjorta, observera flodstranden när de ro längs.
Man håller tre brinnande käppar medan man står nära en lekplats.
Killen håller en svart pinne framför en lekplats.
Två unga flickor leker, den ena bakom den andra.
En ung flicka som gör ett trick mitt i luften framför ett träd.
En man stöttar en pojke när han spelar på en lekplats.
En hund försöker leka med en boll som kastas till den.
Barn i blå koffertar stänker i blå barnpool
Ett litet barn klättrar på en stor vit sovande hund.
En medelålders man i brun hatt iakttar en utomhusmarknad.
Två konståkare, en knäböjande man i svart väst och en kvinna i en skinande gyllene klänning, snurrar ihop på isen.
Den unga pojken i röda jumpos i pölen.
En grupp på 5 barn är klädda i vinterkläder som leker i snön.
En man i jeans ligger på ett trägolv.
En kvinna i en tank topp och en man med lockigt hår spela gitarrer och sjunga i mikrofoner.
En skateboardåkare åker nerför en avsats bredvid trappan.
En man i gul vattentät jacka och hans följeslagare är på en båt i öppet vatten.
Snälla, hjälp min familj här i Kenya.
Två män i täcken gräver ett hål med en spade och några maskiner.
En ung flicka i en blå och grön jacka slädar.
En man och hans söner har kommit till en liten vattendamm.
En flicka som dyker i en allmän pool och njuter av vattnet.
En ung flicka i en grön skjorta som håller en fotbollsboll medan hon står i grönt gräs.
En man med glasögon står framför ett snöigt berg.
En man som bär bast och svarta glasögon slår glatt sönder sin cello på gatorna i ett stadsområde.
Mor och barn går nerför stigen i en lugn takt.
En ung flicka sätter sin fot på marken för att ge balans medan hon cyklar genom parken.
Små barn leker på ett grönt gräsfält.
En tjej med en slingshot i trä, står vid trädgränsen och drar bandet på slingshoten tillbaka.
Ett barn är i luften på en studsande karneval attraktion.
Män klädda i khaki håller en man i armarna.
Män med lövkronor står i ett störtregn.
En mamma som hjälper sin lilla dotter med skidorna en solig dag i backen.
Två män boxas en ring medan en boxare slår den andra.
Två människor ler mot kameran när de åker upp för ett snöigt berg.
En skateboardåkare använder en halv pipa medan folk tittar på.
En pojke med gul hatt och en skjorta som säger "Elmo" pekar mot pannan.
En vuxen och ett barn bär skidutrustning i snön.
Dessa två människor använder årorna för att navigera i havet.
En grupp barn som tränar i ett gym.
En liten pojke som åker skridskor på sin bräda och är redo att slå.
Två män dukar ut den i en boxningsring.
En ung asiatisk flicka glider nerför en stolpe på lekplatsutrustning utomhus.
Musiker mitt i en stor publik.
En liten flicka i gul klänning med röda blommor blåser en vissla.
En liten pojke har pekfingret i munnen.
En man i blå regnjacka som fiskar under en regnstorm.
Ung man åker skridskor på en väg, en solig dag.
En man med isklättrande utrustning klättrar upp på ett istäcke.
En grupp människor står på ett berg i snön.
En ung flicka med långt brunt hår och en röd släde leker i snön.
Olika personer på en brygga med utsikt över havet.
En avliden flicka i en ljusrosa skjorta observeras av en annan flicka i en ljusrosa skjorta.
En bonde som plöjer sin åker med hjälp av två oxar.
En man sitter på en klippa högt uppe i bergen.
En man i grått på en klippa med utsikt över bergen.
En äldre man sitter på en buss och tittar ut över landskapet.
Ett oskyldigt barn utforskar vad naturen har att erbjuda
Två män med orangea skyddsmössor inspekterar stubben i ett nyligen hugget träd.
En ung flicka sitter i gräset och beundrar en liten växt.
Två pojkar försöker äta en banan och ett äpple på soffan, men de distraheras av förvåning.
En tjej sitter på en killes knä på en fest.
En kvinna i orange arbetskläder bredvid en stor blå soptunna hjälper en man sopa lite smuts och vatten i en soptunna.
En man sveper ut medan han bär ett barn på ryggen i en hållare.
En kroppsmodifierare njuter av en öl samtidigt som den slappnar av på en trevlig solig dag.
DJ-killar som är dumma för kameran.
Ett marschband övar på ett utomhusfält.
En skäggig man med brun skjorta spelar gitarr.
Barn spelar 3 på 3 pingis i ett gym.
Två män spelar en dubbel tennis match.
En röd racerbil med en förare i en himmelsblå hjälm i racingbanan.
En person med svart jacka hoppar i snön.
En ung flicka med långt svart hår klättrar på en bit rep lekplats utrustning.
En man och en kvinna sätter sig i boxningsställning för att börja träna.
En grupp dansare, som bär svarta byxor, tanktoppar och svarta hattar, dansar och håller käppar i luften, med sina högra ben något utsträckta.
En man som håller i en mikrofon och täcker ögonen
En familj som håller händerna i snön är bakom en man och hans son, som bär en blå jacka.
Två flickor med anka som flyter hoppar ner i mörkt vatten.
En kvinna i grå klänning och höga klackar som håller ett barn i rosa klänning medan hon stirrar ut en glasskjutdörr.
Människan identifierar trädslag för unga par under snöskovandringen.
En asiatisk flicka som bär en Camelbak och går skor och går sin hund i en snöig skog.
Två unga pojkar bowlar med stötfångare.
En joggare med en hund som springer mot en brandbil med förlängd stege på en väg
Två damer som joggar på en stig nära vattnet.
En ung pojke vid 13 års ålder leker i snön och har en snösko på benet, och springer
På det här fotot blir män hedrade för sitt mod.
En pojke i orange jacka klättrar genom en lektunnel
En kvinna som lagar mat över en öppen härd.
En grupp afrikanska barn visar symboler skrivna på krittavlor mitt i ett smutsfält.
En pojke sparkar en boll i sitt vardagsrum.
En man har klättrat upp till toppen av en röd ljusstav och rör vid ljuset.
En skateboardare utför tricks på ett hopp från en ramp.
En ung kvinna i svart blus läser en bok på ett plan.
Pojke i röd skjorta stående på taket av en byggnad medan ett annat barn tittar på underifrån.
En person som bär en mörkblå mörkklädd klädsel från huvud till tå, med mask och väst och håller ett tunt svärd.
Några män spelar volleyboll.
Labbet tittar genom ett mikroskop i ett labb.
Q barn i röd skjorta skapar en rock utställning.
Tre äldre kvinnor stannar för att titta på en utställning i ett museum.
En vetenskapsman tittar i sitt mikroskop.
En ung dam rider en brun och vit häst.
Publiken tittar på färgglada varmluftsballonger i fjärran.
En liten pojke använder ett teleskop för att se ett objekt långt borta medan en liten flicka står i närheten och tittar.
Människan håller en linje när varmluftsballongen är uppblåst.
Stora grupper av familjer samlas på en utomhusgård för att be om regn.
Den lilla pojken bär vita shorts.
En snowboardåkare med röd rock går nerför en snötäckt sluttning.
En kvinna som har en blacker top dans framför ett band.
En grupp unga vuxna är organiserade en varm dag i en park med en fontän.
En man med skägg, rött pannband och läderväst ler.
En pojke hoppar in i en pool och visar ett fredstecken till kameran.
En kvinna i en handduk slappnar av i en bastu.
En kvinna med en väska står på en gata nära en man som lutar sig mot en vägg.
Cowboy håller i hästen
Två kirurger arbetar hårt med att undersöka en patient.
En manlig tonåring rider nerför en snötäckt kulle i en grön släde.
En skidåkare lutar sig åt ena sidan för att gräva sina skidor i snön.
Män förbereder sig för att skjuta med sina vapen.
En ung pojke i en långärmad t-shirt tittar upp på kameran från ett öppet område långt över marknivå.
Man sitter på en gammaldags vagn.
En monsterbil flyger genom luften framför en arena fylld med åskådare.
En man har smink applicerat på sitt ansikte.
Tangentbordisten och en kvinnlig sångare delar en mikrofon medan en andra man tittar på.
En man utan tröja som jobbar på ett tak.
Det finns en man som arbetar på taket av ett hus som antingen håller på att nybyggas eller byggas om.
En skjortlös man som bär blå jeans går längs ett gräsigt område.
En tjej i grön skjorta spelar på en gunga.
En man hugger upp mat på marken.
Två munkar i traditionella apelsindräkter går nerför en trappa.
En skjortlös, handskebyggd byggnadsarbetare står på ett skenat tak.
Det finns flera personer men i synnerhet tre, kommer från ett köpcentrum med lådor och växter i sina vagnar.
Ett litet barn, nappare i munnen, står med händerna upp mot en glasdörr och tittar ut.
En jordgubbshårig kille blinkar med sina blå ögon och ett stort leende mot kameran.
Två flickor sitter vid en dörröppning på trappan.
En pilot sätter sitt bagage bredvid planet på flygplatsen.
En publik tittar på många på en cykel utför ett stunt.
Två män på en blå kanot mitt i en stor vattensamling.
En kvinna i jeans klättring.
En manlig dansare i beige lyfter upp sin kvinnliga kamrat på axeln, när hon svävar över folkmassan.
Två indiska kvinnor sitter på en marknad bakom grönsaker.
Person med skidstav och röd jacka, går på ett snötäckt träd över vatten.
En far med 3 barn tittar på en målning av en skogbevuxen bergsscen.
En asiatisk kvinna, och en svart man, går förbi trapporna till tunnelbanan.
En man håller på att ramla ner från en stege.
Tre kvinnor och två män använder triangelformade nät i en ström.
En vandrare utgör för en bild framför fantastiska berg och moln.
En ung kvinna gör uppskjutningar framför tre medlemmar av de väpnade styrkorna vid ett konferensevenemang.
En ung vuxen ler efter att ha glidit nerför en snöig, nedsänkt kulle.
En liten pojke med en orange jacka gräver i sanden bredvid en flagga.
Tre män och en pojke rider en orange berg-och dalbana.
Poliser i upploppsdräkt, tillsammans med två poliser på hästryggen, anklagar en folkmassa som är bakom en barriär.
Två barn, en i vit skjorta och en i svart skjorta, liggande på kuddar.
En dansare i en rosa tutu slår en pose utanför en byggnad som är täckt med graffiti.
Tre små barn på en sten, tittar på vattnet.
En grupp indiska unga kvinnor och flickor badar vid kanten av en pool med sina torra kläder och en byggnad i bakgrunden.
En blond kille i grön tröja äter en smörgås.
Den här lilla flickan, hennes blonda hår hålls tillbaka av ett rött band, sticker ut tungan lekfullt vid kameran.
Några unga flickor i ett klassrum.
Kvinnan slappnar av genom att doppa fötterna i vatten i ett stenigt område.
Flera män i svart och vit rutig duk, dansar runt en fackla.
En man med orange skjorta plockar upp en fritös med ätpinnar.
En kvinna med lila skjorta i solglasögon, liggande på sin bokväska.
En kvinna i en ljusrosa tröja som kastar en fiskelina i en sjö.
Tröjlösa män i matchande kläder lyfter händerna upp i luften.
Skateboardaren i en vit t-shirt och blå mössa sitter på sin bräda och kustar ner i den milda klass.
En man sitter på en skateboard på trottoaren.
En basketspelare i vit uniform försöker blockera ett skott från en basketspelare i en mörkblå uniform.
En kvinna handlar färsk mat på en utomhusmarknad.
En grupp barn sitter nära varandra och skrattar medan en pojke i vit skjorta hoppar över dem.
En kvinna sitter vid ett teleskop.
En ung kvinna klädd i lila kostym med vita vingar ger en liten pojke i en blå jacka en bit godis.
En boxare försöker slå sin försvarsmotståndare med ett våldsamt uttryck i ansiktet.
En vandrare i snöskor ute för en promenad i snön pauser för att titta på kameran.
Ungdomar joggar i snön i den här stadsscenen.
Mina herrar med en svart och gul skjorta står på scenen och spelar gitarr.
En grupp människor vandrar genom isen.
Unga människor på skateboard och en utan tröja hoppar i luften.
En grupp människor skrattar med böcker i bakgrunden.
Två anställda knådade och förbereda deg för användning med att göra kakor som syns genom fönstret.
En kock i vita kläder sätter något i en tegelugn.
Två män som verkar vara matförsäljare kör en röd kärra full av frukt.
En man går genom ett fält med något slags trädgårdsredskap.
En man hukar sig på sin åker och skördar rötter mitt på dagen.
Två män i en fält eller djungel tittar på något.
En person som snowboardar nerför ett berg täckt med färsk pulver snö med tallar i bakgrunden.
En skateboardåkare på en skatepark som försöker sig på ett järnvägsspår.
En man i en röd jacka använder en maskin på isblock framför flera åskådare.
En liten vit pojke klädd i vinterkläder stående vid ett träd i snön.
Flera personer arbetar i den varma tillverkningsanläggningen.
Skidåkare som snöas på när de korsar snölandskapet.
En man i vit skjorta ler när han säljer sin gatumat.
En ung person slädar nerför en kulle i snön.
Person som bär en lila rock sittande i snön under ett träd och äter en smörgås.
En man som skulpterar en liten lerkruka på ett spinnhjul
En man i vit skjorta och jeans sopar trottoaren på en gata.
En asiatisk dam står med en vagn med potatis.
Påven och en annan man i svart kostym har ett samtal.
Ett barn utan tröja som springer i smutsen.
Flera höga kvinnor hoppar upp i luften samtidigt bär traditionella matchade kläder och sandaler med tre alfta varmluftsballonger i bakgrunden.
Barn arbetar på ett uppdrag i skolan.
En man och en kvinna dansar tillsammans.
En liten flicka håller en snögubbes grenade arm.
En skäggig man med blå randiga shorts, en mörk tee-shirt och baklänges baseball keps står vid ratten på ett fartyg som flyger en söndersliten röd flagga öppet vatten.
En man är på en båt på lugnt vatten och har repet.
Små barn i röd jacka och khaki byxor på toppen av en rutschkana med ett staket bakom.
Det finns flera människor utanför som tittar på ekollon squash.
En flicka som knäböjer i vad som verkar vara en kyrka.
En man böjer sig bakåt med svarta remmar runt sig.
Silhuetten av en person som hoppar i luften under en solnedgång.
En man som väntar på att trafiken ska stanna vid vägkorsningen
En gul slang sträcker sig från en av två benvita fordon parkerade bakom utsträckta försiktighetstejp, som flera figurer samlas på trottoaren.
Brandbilar och andra nödfordon reagerar på en nödsituation.
En man i en traktor som kör på en dammig väg!
En präst i telefon nära några kvinnliga militärarbetare som tar en paus.
Börjar en omgång hårhockey mellan två män.
Två kvinnor och ett barn som sitter vid en sten med stickade saker.
En grupp asiatiska människor som tittar på hantverksmateriel som erbjuds av en ung kvinna.
Två barnsläde som rider nerför en kulle.
En brandman är på taket av huset.
En ung person tittar blygt på kameran.
En ung pojke i röd dräkt som håller en skotrofé ovanför huvudet.
En person i en rock läser en tidning på en bänk.
En barfota man i svarta shorts sover på en dörr framför en röd dörr.
En nyfödd med en skjorta som säger: "Jag är chefen."
Barn deltar i ett säcklopp utomhus med många andra barn som observerar i närheten.
En pojke sjunger in i en mikrofon, scenljus i bakgrunden.
En man som hoppar från en dykbräda till en pool.
En gymnast snurrar ett vackert band.
Ett barn som bär blå skjorta och shorts gräver ett hål i sanden nästa två en liten grön spade.
En ung brunett flicka bär en Toronto Maple Leaf skjorta poserar med en hockey pinne och puck.
Ett spel av rugby där 2 spelare försöker stoppa det motståndare från att fånga en boll i luften.
En pojke i orange skjorta sitter på en sten nära vattnet.
Ett ungt barn gråter medan han eller hon knäpper sin pyjamas.
På fiskmarknaden mäter en arbetare och filar en fisk.
Många arbetare med blå skjortor och vita förkläden förbereder fisk till salu.
En professor i svart blazer är författare på en krittavla.
En grupp unga män står och sitter runt en brandgrop medan de dricker och grillar sin mat.
En liten flicka i ett vitt badkar håller ett träföremål i vattnet.
Ett fordon som bär hö rymmer också en ung pojke och två män som sitter ovanpå höet.
Två personer gömmer sig under jätteskålar, kanske för att undvika solen.
Det finns en äldre man som stryker en skjorta för sitt arbete.
Flera pojkar leker ute på fältet.
Två unga flickor rider en stor cykel på sidan av vägen.
En liten pojke som leker med en pistol.
En man skriver något på en markörtavla i ett klassrum när någon tittar på honom.
Två män brottas på mattan medan publiken tittar på.
En vit man med svart hår klädd fint i grå klänning byxor, blazer och lila slips står på gatan framför ett garage vända en pannkaka som fångas i luften.
En ung pojke och 2 flickor öppnar julklappar.
Ett ungt rödhårigt barn är på väg att ta en tugga av ett blått fruset mellanmål.
Sex barn sitter runt ett rektangulärt matbord med en grön duk och mat på.
Två flickor ligger mag-ner i gräset samtidigt dela hörlurar till en mp3 spelare.
Två flickor lutar sig bakåt på däck gungor och ser upp och ner på kameran.
Två män står i en lyftkran bredvid flera höga träd.
Cowboy börjar ramla av en knocking bronco.
En person visas upp och ner på sin cykel över ett stort fält.
En cyklist gör ett stunt medan åskådare tittar i det avlägsna hörnet.
En kvinna går över en stege mellan två berg.
En kvinna i svartvitt som korsar en väg.
Två äldre kvinnor handlar blommor medan en afrikan-amerikan man tittar på deras sida.
Två barn leker i nuet och rullar in det i en stor boll.
En ung blond pojke tittar på en röd hundskål och en sjaskig hund sitter bakom honom.
Två pojkar som använder krita för att skriva på trottoaren.
Ett barn i vit skjorta är nedsänkt i en sving framför tvättmaskinen.
En kvinna och en ung flicka rider glatt på en karusell.
Två barn sover i en barnvagn på trottoaren.
Två barn leker läkare med ett spädbarn.
En ung blondhårig pojke åker ner för en röd rutschkana.
3 man spelar musik tillsammans bestående av gitarr, violin och banjo.
En äldre man i en blå skjorta som står mot en svart pipa.
Fyra poliser patrullerar på gatorna på hästryggen.
En man med solbränd hatt och skjorta, en orange skyddsväst och mörka glasögon gester mot en närliggande bil.
Långhårig man jobbar i ett vitt rum.
En man med en svart jacka spelar på sin smartphone, medan den lilla flickan bredvid honom bär en scarf och blå jacka läser en bok.
En man ska fiska på sin båt som kallas Melanie.
En dam ler medan hon sitter framför hela maten och håller ett matobjekt.
En tjej i röd skjorta är i en bowlinghall.
En besättning gör ett plan redo att lyfta.
En tunn medelålders man står bakom ett podi i ett tomt bankettrum.
En snowboardåkare fångar lite luft från ett hopp på ett snötäckt berg.
En äldre gentleman med ansiktsfärg spelar fiol.
En ung pojke kysser en man i pannan när han sover.
En man som står framför flera jordhögar om spade med andra.
En soldat klädd i stridsredskap skalar en mur för att förena sig med sina kamrater på andra sidan.
En man inspekterar skador i ett förstört rum.
Det finns en man som bär svart och vitt sittande på en stolpe med deras ansikte målade vita håller bollar.
En pojke tar något från en låda som hålls av en man i en kanin kostym.
Ett blond barn som sover i sängen med en filt ovanpå sig.
En person som använder en stege för att måla en kolumn vit.
En man i vit skjorta och grön väst använder gamla verktyg för att forma en bit trädstam.
En byggnadsman med blå hatt stirrar ner under.
Två arbetare i hårda hattar och säkerhetsselar reparerar ett tak.
En ung man är på sin dator i en kontorsmiljö.
Två kvinnor bär förkläden och bakar kläder och lagar något i ett kök.
Två pojkar fick stryk bakom ett hus och lämnade det.
En man arbetar i en konststudio och är omgiven av konstartiklar.
En liten flicka som skrattar medan hon går ner i en rutschkana.
Tjejen sitter på en stol och sms:ar på sin telefon.
Jag ser en grupp människor stå runt omkring och en polis stå runt.
Mannen är stolt över sitt hantverk när han koncentrerar sig på sin snidning.
En dam med en röd väska lämnar affären.
En skäggig man och en blond kvinna sitter i publiken
Hårdhackade byggnadsarbetare väntar på att få gå ombord på en hiss.
En man äter mat på ett bord framför en liten mataffär på gatan medan en förbipasserande går förbi.
En kvinna i lila kysser ett barn efter hennes uppträdande.
De lokala barnen har en fotkapplöpning.
En tjej i vit skjorta springer.
En klättrare stannar för att ta en drink medan han klättrar på ett snötäckt berg.
En man sitter på en snöbank.
Två barn leker i en utomhuspool.
Två män på en parkeringsplats i ett företag en man tittar på den andra mannen hoppa.
En musiker som spelar en scen upplyst i rött sjunger in i en mikrofon.
En person är upp och ner och gör en volt på en snowboard.
En man sitter på en stol framför en hög vattenmeloner.
Fyra dansare i gult framför en etnisk dans.
En man i blå snödräkt gör en volt på ett stort snöigt berg.
En fiskare skär bete ombord sin båt, som är förtöjd vid kajen, medan pelikaner simmar i närheten.
En äldre metallarbetare slipar ner en bit plåt i en verkstad.
En man på en cykel leder en annan cykel längs en stadsgränd.
Två barn, hopslagna mot kylan, byggde en liten snögubbe.
Tre män sitter och funderar på sin nästa tjurtur.
Ung man, i sönderslitna byxor, sitter på avsatsen i ett fönster och spelar fiol.
En kvinna blandar ihop en smet av mat.
En grupp svarta barn poserar för kameran.
En köpman poserar i en slaktarbutik.
Två pojkar kanonkulor i en sjö nära en röd paddelbåt.
En man som sitter på sin arbetsplats och gör smycken.
En indisk man arbetar på en textil i bakgrunden medan en indisk kvinna arbetar med färgämnen i förgrunden.
En parad av folk som bär röd marsch förbi en byggnad medan de spelar instrument.
En man hukar sig ner medan han målar sina konstverk på en stor garagedörr i metall.
Flicka som utför ett hopp i luften med hjälp av ett sidenband.
En pojke med röda solade skor leker på en gunga.
En vithårig gammal dam, klädd i en rutig skjorta och shoppat.
En ung kvinnlig gymnast ligger ner på en matta medan han tittar på en hula-hoop.
Ett kamerateam förbereder sig för att filma med en videokamera.
En nyhetsutgivare i en blå rock ger sin rapport i regnet.
En ung man fångar lite luft medan han rider på en vågbräda.
En man i blå jacka knäböjer på en strandpromenad bredvid havet så att han kan justera sin fiskespölina.
Person i motion kläder klättrar ett rep.
En man utövar all sin kraft i ett gym med en stor mängd tyngdlyft över huvudet.
En trafikpolis leder trafiken i ett stort befolkningsområde.
En pilot med hörlurar sitter i sittbrunnen med sin andrepilot.
Ett barn som leker med stenar.
Grå hund kör ner trottoaren mot tvättlinje på gårdsplanen.
Två personer som sitter nära en dörr och håller skålar i knäna.
Tjejen leker i en pöl med bara fötter.
En man klär sig i sitt hem när han tittar på sin laptop.
Ett barn som sitter på marken, ser ut som hon är djupt i tankarna.
En tonårspojke och en flicka som njuter av fondue.
Två män, en i blått och en i rött, spelar hockey på ett plan.
En dam i en zebra-strippad rock interagerar med någon klädd i en pandadräkt.
En grupp unga pojkar spelar baseboll i ett främmande land
Tre män jobbar med sina cyklar i axeln på en väg.
Kunder och arbetare vid kassan i en butik med röda diskar och kundvagnar.
Två män som bär svarta skjortor och byxor håller i träpinnar.
En man i beigedräkt spelar trumpet i en mikrofon.
Tre kvinnor deltar i en dans på en campingplats.
En livemusikkonsert släpper konfetti från taket medan publiken hejar på, exstatiskt.
En kvinna som hoppar framför en graffitivägg.
En ung man sträcker på benet och balanserar en skiva på fingret.
En grupp studenter som spelar Jenga.
Två asiatiska kvinnor sitter i ett gathörn, medan en vit bil passerar förbi.
En stor flicka med blå jeans hoppar över en stubbe.
En man som arbetar på fälten när han rör händerna runt det höga gräset.
En ung dam tar sig tid att tänka på en offentlig bänk.
En kvinna klädd i cosplay utanför visar upp sig för kameran.
En kvinna i snöskor tittar på ett papper.
En hand håller en penna över en sida med noter.
En kvinna i en godisaffär som surfar på godis.
En kvinna tittar in i en soptunna utanför Mango Mang.
En dam lagar en annan dams hår.
En äldre man i orange skjorta och gröna shorts går förbi en byggnad dekorerad med graffiti.
Två barn spelar fotboll på grönt gräs.
Fiskare på båten tar tag i ett nät fyllt med vad som verkar vara musslor.
Confetti är i luften bland en stor skara människor vid någon form av firande.
En sångare är het och svettig från att uppträda i en konsert.
Polisen tittar på varandra på hästar.
En man som håller ett barn tittar på leksaker i en affär.
En fotbollsspelare sparkar en boll.
En kvinna i svart skjorta, med en halsduk runt halsen, syr.
En polis med många föremål runt midjan beställer något på ett café.
En färgglad målad och klädd man uppträder för publiken.
En kvinna som knuffar en kundvagn i en mataffär.
En man som bär solglasögon sitter i ett vitt fordon med ett vapen på dörren.
En pojke ler omgiven av flera andra människor ler mot kameran.
En man med glas och en kvinna med rosa skjorta sitter bredvid varandra.
En man talar på ett podi i en kyrka.
En kvinna med handen i en stor kruka vid en vattenpump utanför.
Två vuxna kvinnor, en med paraply, och en liten flicka som går på en bro.
Flera personer, däribland en kvinna i röd klänning som håller ett barn, befinner sig på en gata nära dussintals duvor.
Ett litet barn hänger ut genom fönstret på en buss.
Fyra män i lila skjortor och två i mörkgrå med en skulptur.
Människor som arbetar tillsammans fyller skottkärror på en lekplats.
En grupp unga fotbollsspelare springer nerför planen efter bollen.
En skidåkare flyger genom luften medan han gör ett trick.
En manlig surfare som föll av sin surfbräda ovanpå en liten våg
En äldre man och en ung flicka tittar på fisken i en konstgjord damm.
En artist knäböjer vid kanten av en scen för att få något från en kvinna i första raden.
Två män hoppar från marken under en sparring tävling mellan motståndare.
Ett äldre par dansar bredvid ett bord där en pojke sitter med huvudet nedåt.
En ung kvinna, som bär på flera väskor, hoppar upp i luften.
Två kvinnor bär röda etniska dräkter, med en kinesisk byggnad och ett berg i bakgrunden.
En man och en pojke som rör varandras händer med två andra människor i bakgrunden.
Två män simmar på en strand med en trädtäckt kulle i bakgrunden.
Pojken spelar volleyboll på stranden.
Två män spelar boll, en vit en svart, med den svarta hoppar mot höger sida av ramen.
Sju personer använder PC-bord i ett rundat bord.
En man i grön jacka har satt upp en kamera på några stenar.
En man som står framför en träbro nära en stenig flod.
En man med nyanser och en svart skjorta på att uppträda passionerat på scen.
En grupp barn njuter av snacks och spelar ett brädspel tillsammans.
En forskare i ett labb pekar på en datorskärm medan en av hans medarbetare tittar på.
En snowboardåkare i luften med ljusgula byxor.
En byggnadsman tar en paus medan han tittar på utsikten.
En stadsgata har tre personer som går i olika riktningar.
En man klädd i en traditionell infödd amerikansk klädsel spelar ett instrument infödda till sitt folk.
En kvinna i brun klänning hoppar från några trappor utanför en byggnad.
Vissa anställda i gula skjortor hjälper till med lokala barn i konst och hantverk.
En man, med en röd sporttröja, tittar på en fotbollsmatch.
Fyra killar i vita labbrockar med skåp i bakgrunden som håller något i brand.
En kvinna i rutig kjol och en man med rutiga strumpor, kilt gör sig redo att dansa natten bort.
Flera människor som ligger ner på en stenig strand i förgrunden med människor som står upp i bakgrunden.
En grupp människor dansar i färgglada kostymer framför en Fired Earth-butik.
En grupp kvinnor, klädda i festliga blå klänningar och fjäder huvud inredning, parad nerför gatan.
Två kvinnor som spelar framför en dörr märkt "The Castle Keep".
Tre unga damer i gul uniform tar en paus vid ett litet bord.
En man i svart hatt och shorts kastar en matchande gul glöd pinne
En ung dam med vild blont hår spelar elgitarr på scenen.
Fyra barn leker i sanden nära vattenbrynet.
En fotbollsspelare i röd uniform är på väg att sparka bollen.
En liten flicka borstar tänderna.
En skara åskådare på en traktortur ser på när en jordbrukare arbetar hårt ute på fältet.
En man med en kundvagn studerar hyllorna i en snabbköpsgång.
En man står på byggnadsställningar i en studio medan en eld brinner i förgrunden.
Ett actionfoto på scenen i ett punkrockband.
Ett par, som såg ut som Aladdin och Jasmine, rider den magiska mattan på en natthimle.
En svart och en vit hund jagar en tennisboll.
Glada, leende småbarn sitter i en ganska blå, vit och gul filt kasta en stor blå boll.
Ett band framför en låt på en klubb.
En ung pojke som håller andan och hoppar i sjön en varm dag.
En grupp kvinnor i saris sitter, pratar och badar tillsammans.
En pojke i vadderad hjälm studsar på en studsmatta inomhus.
Den här arbetaren kör sin vagn genom den livliga trafiken ensam.
En gitarrist jams för en publik på hans röda instrument omgiven av hans band kompisar under strömmande vitt ljus.
En man spelar dragspel längs gatorna, underhållande förbipasserande.
En skara vuxna som är klädda i ljusa färger klappar händerna.
En tjej spelar fiol och en klarinett bakom sig.
En kvinna i randig skjorta går en häst tvärs över en gata.
En man observerar en målning medan en annan person försöker återskapa samma målning.
En motorcykelpolis undersöker en ljus neonreflekterande väst medan han står bredvid två färgstarka polis motorcyklar.
Ett litet barn leker med leksaker i en träbänk.
En man i ett vitt förkläde grillar på en grill utanför.
Fyra män hänger på möbler medan alla sitter på sina bärbara datorer mot en solbränd vägg.
Det finns en man i en röd tröja som försöker göra ett trick på en skateboard.
Flera människor i kostymer från Disney-filmer går nerför en gata.
En turnégrupp sitter på den andra historien om en dubbeldäckare turnébuss mitt på Times Square.
En vacker dam sitter ner och öppnar sin väska.
En man som åker vattenskidor med vattnet som flyger upp bakom honom.
En äldre kvinna som rullar ut deg att baka med.
En man som är delvis skallig med solglasögon på, en svart tröja och jeans, har en spade och skyfflar trottoaren och några trappor medan en gyllene retriever tittar på honom.
En man och hans kvinnliga assistent använder en propanbrännare för att grilla biffar.
En person som plockar garbanzobönor med sina björnhänder.
En man färdas med två åsnor i bergen
En ensam klättrare på ett snötäckt berg med flera stora berg i bakgrunden.
En skäggig man i blå jeans på en skateboard hoppar över en kundvagn.
Två personer klättrar genom ett nät av metallsträckor med shorts och tennisskor.
En man maler ner en räls på en skateboard.
En kvinna med ljusa röda läppar och en randig skjorta är ansträngande framför en mikrofon på ett stativ, medan en annan person är i bakgrunden håller en mikrofon.
En ung pojke lagar kött på en grill utanför.
En asiatisk man, kvinna och pojke väljer paketerad mat på en innermarknad.
Ett marschband med blå och svarta danser på gatan.
Två barn står och möter kameran framför ett dinosaurieskelett.
Två personer, en man och en kvinna, hoppar samtidigt.
En ung flicka i karateuniform hoppar från en studsmatta när hennes instruktör ser på.
En tjej som bär rosa hänger på korgarna.
Ett barn, som sitter vid ett bord med kritor och konstartiklar, ritar en bild med ett barn i bakgrunden.
En kvinna med mikrofon som gör espresso
Någon i en regnjacka skjuter en gul väska på hjul nerför trottoaren.
Små pojkar som spelar fotboll bär orange och svart
Ett lag av pojkar i röda och svarta uniformer spelar fotboll på en plan.
2 asiatiska män sveper blomblad från några trappor.
En person i svarta pannor och en svart t-shirt hoppar på en fontän plaza.
En grupp pojkar bygger något med trä.
Två kvinnor skyfflar jord på en gård vid ett stängsel.
En man som bär skyddsglasögon reparerar ett cykeldäck.
En man i svart utstyrsel, med lågor på, övar sin kampteknik.
Barnet går genom högt gräs en solig dag.
En flicka verkar hänga upp och ner från ett djungelgym.
En unge upphängd i luften av några kablar.
En idrottsman i röda shorts fångas frusen under ett basket drag.
Flickorna återvänder till fältet under sin softball match.
Två män i skeppet "Amble" ställer ut lastade med fällor.
Två hundar springer i smutsen
En kvinna som bär en svart och blå klänning figur skridskor på ett ben.
En liten pojke tittar på sitt teleskop på dagtid.
En äldre man med vitt hår och skägg pratar in i en mikrofon.
Byggarbetare använder kablar för att hänga från byggnadernas sidor.
Två små flickor står på en liten avsats med sina ansikten mot en tegelvägg.
En pojke som håller i en skateboard hoppar över en annan pojke.
En man och en kvinna klädda som motorvägsanställda jobbar på sidan av vägen.
Flera statliga arbetare som arbetar på en järnvägskorsning.
Färgfullt klädd man dansar på gatorna, samtidigt balanserar något på huvudet.
En kille som snowboardar nerför ett stort berg.
En skidåkare åker skidor nerför ett berg med goggles och en röd anorak.
En man är på sin mountainbike och flyger i luften.
En man sitter och säljer blommor och grönsaker på en livlig gata.
En person som går med sin cykel och två andra människor.
En man med skägg reparerar ett nät som sitter med en boj och rep bredvid honom.
En person kommer in i baksätet på en lastbil medan arbetarna arbetar bakom.
En man med ett hårigt bröst klipper en gräsmatta.
En pojke med randig skjorta sitter vid ett bord och skär något.
En leende pojke gör en gest med ena handen samtidigt som han håller en stor flaska läsk i den andra.
Ett barn och en kvinna utför trädgårdsarbete.
En man som hoppar sin cykel från jordhögar är flera meter i luften.
En terrängcyklist rider över en stock.
En man på gatan spelar sin gitarr för publiken.
Två kvinnor handlar mat i affären.
En kvinna väntar med barn när hon checkas ut på Walmart.
En äldre man handlar tvätttvål på Walmart.
En kvinna i bikini står i vatten och är omgiven av fisk.
Två män utan skjortor är på taket.
En äldre man i vit skjorta tittar på en webbsida på sin dator, på sitt kontor.
Officeren på den vita mopeden går över kullerstenspromenaden.
En man på en cykel rider förbi en gul byggnad som har markerats med graffiti.
Kvinna sätter upp ett fotografi av en gentleman i rullstol med 3 åskådare och två tjänstemän.
En man klädd som kolonist talar till en folkmassa i en molnig stad.
En man som leder en orkester och undervisar människor.
En man med en kamera på axeln videofilmar en konsertuppvisning.
Man klipper gräs nära en byggnad med ansiktskläder för skydd.
En man är ute och tvättar sin bil med tvål och vatten.
En kvinna utför gymnastik med långa röda band.
En kvinna i solglasögon som gör ett surande ansikte medan hon äter skaldjur.
En man i neonkläder fixar en gatuskylt.
En medelålders kvinna sopar trottoaren framför en butik i en stad.
En man som städar fönstret i en presentbutik.
En man i uniform sitter på en ramp och tittar tillbaka på en staplad rad matvagnar.
Damerna i lila jackor spelar sax.
En grupp män i shorts och skjortor som joggar längs en tegelgång.
En grupp män står vid en vit lastbil.
En man torkar upp insidan av en nöjespark rida som är täckt med blå plastlakan.
En man kör en vagn på en gångbana.
En manlig gitarrist sjunger kraftigt en inte till en låt i ett dåligt upplyst rum.
En man som spelar dragspel med en flicka som sjunger och spelar tamburin.
En förväntansfull kvinna låter glatt en annan lyssna på barnet inuti henne.
Två personer knuffar en kundvagn på en folk-mover.
Två män sitter i en fortkörningsbåt i vattnet, med land- och segelbåtar i bakgrunden.
Två uniformerade män rider i en motoriserad båt.
Flera män i flytvästar och andra redskap på en båt i vattnet.
Bandet med fyra killar uppträder på en ljust upplyst scen.
Fem kvinnor, som bär långa infödingsdräkter, och två män, som bara bär byxor, visas i vattnet, samtalar och plaskar.
Man klädd upp är färgglada kläder gör ballong konst.
Två personer som tävlar med lansar och sköldar på hästar medan människor vaktar från under ett tält och utanför tältet.
En man i hjälm rider en ATV i en öken.
En ung flicka med polka prick klänning och kanin öron spelar ett arkadspel.
En man torkar utsidan av ett fönster rent som en flicka rengör samma fönster från insidan.
En man med vit t-shirt och blå jeans gör ett handstånd på en grön gräsmatta.
Två män tar bort trädgrenar.
Tre kvinnor i klänningar står på en scen och lutar sig tillbaka på ett ben med en gardin bakom sig.
En grupp unga vuxna som hejar i en folkmassa.
En plattform flyter på en flod med en man som spelar piano, en kvinna som sjunger och en man med åra roddar på plattformen.
En man som drar en rickshaw eller handvagn delar en väg i Kina med en Audi och lastbil.
Fyra män försöker fixa en varmluftsballong med en annan varmluftsballong sedd i bakgrunden.
En man rullar på ett räcke.
En ung man glider nerför en ledstång på rullskridskor medan folk bakom honom tittar på honom i parken.
Flera brandmän står utomhus i full uniform
En man i en klargrön skjorta och hård hatt klättrar upp i ett träd.
Vägarbetare bär orangefärg på en arbetsplats.
En liten flicka borstar tänderna med en orange och blå tandborste.
En hane med solglasögon petar på ett träd med en stolpe.
Två män som använder en slang som hänger ner i vattnet, målet för den är oklart i bilden.
En grupp människor i uppblåsbara flottar som försöker manövrera i en isig flod.
En liten flicka i en flytväst i havet tittar på en val bredvid båten.
Underhållsarbetare som städar sidan av ett rött och vitt tåg.
En gammal man i blå skjorta cyklar förbi ett stort kryssningsfartyg.
Kvinnan arbetar med sin symaskin.
En kvinna med blont hår, med ljusa röda ränder på toppen som arbetar på en dator.
Barn leker utomhus i en fontän.
Den unga damen som bär ytterkläder kastar en blå fotboll, med ett par andra människor på fotot som ser ut som studenter, en solig dag.
En vägarbetare i grönt, det finns en orange kon nära honom.
Byggarbetare i blå byxor och limegröna skjortor skar grenar från ett träd.
Tre landskap arbetar bort en fallen trädgren.
En ung blond kvinna i idrottskläder ska kasta en blå fotboll.
En kvinna i svart som ligger på en matta i ett lugnt rum.
Två barn som spelar i en fotbollsmatch på en fotbollsplan.
En tjurryttare, i full stoppning och med hjälm, rider en stor brun och vit tjur.
Två unga pojkar sitter i lådor i vardagsrummet nära några dekorativa stolar.
En kvinna i en ljusröd klänning står utanför en byggnad.
En ung man sjunger på scenen med mikrofonen i munnen.
Ett band uppträder på en liten scen med neonljus som lyser.
En man i neonskjorta, khakis, och en orange hård hatt går förbi en mulchmaskin.
En ung latinamerikansk pojke som sitter baklänges på en åsna.
Familjen sitter på ett gräsfält medan andra går förbi.
En man i en byggnadsdräkt arbetar på att putsa trädgrenar.
En flicka i en grå tank topp ger ett glas till en man i en vit skjorta.
Ett team kockar arbetar för att förbereda en måltid.
En man som bär en hård hatt matar en borste till en industriell flishuggare.
En äldre man håller i armarna på en ung pojke som bär batmanbyxor.
En pojke i en röd jersey spelar ishokey på en utomhusis rink.
Två män, en i svart rock, har ett samtal framför en byggnad.
Två kvinnor med vita huvudskydd stirrar på en mobiltelefon.
Kvinnor pekar ut hennes arm medan hon står i en position.
En man och två pojkar står och sprutar vatten.
Folk går omkring utomhus antingen under höst- eller vintersäsongen.
En äldre kvinna i ett tält använder sax och stol för att reparera ett fiskenät.
De äldre herrarna förklarar med entusiasm vad strängen är till för.
En grupp män som bär cowboyhattar sitter bredvid en häst.
Damen i en ganska ljusgul klänning blir ombedd att dansa, medan barnen ser på.
En kvinna som bär en grön och rosa klänning dansar med någon som bär en blå topp med vita byxor.
En grupp ungdomar som är på väg att uppträda inför en åhörarskara.
Två små flickor i en affär som tittar på barbie leksaker.
En man i vit skjorta står på ett flygplan.
Två män i baseballuniform spelar baseball, en ligger på marken med hjälm och den andra hukar.
Två kvinnliga cowgirls sitter på väl underhållna hästar bär vita hattar.
En man i vit uniform med blå trim tillagar mat för servering.
Två kanoter som flyter nerför floden med varor.
En ung man solar på en vacker strand med ett torn mitt i havet.
Tre små barn observerar och interagerar med ett mikroskop och en dator.
Den här unga kvinnan får manikyr på en salong.
Två män och fyra barn i matchande kläder.
Det är många barn som går på tågspår omgivna av träd.
2 män brottas och är i luften, medan domaren och åskådare observerar.
Här är en bild på en lärare som pratar på en mikrofon i sitt klassrum.
En man på en cykel pratar med en kvinna som sitter bakom några bord.
En tunnelbanestation där många människor står och en kvinna sitter och läser.
Två officerare på hästryggen tittar nerför stadsgatan.
Tränare för North Side baseball laget prata med sina spelare i utgrävningen.
Välklädd man och kvinna dansar på gatan
Denna mor och hennes dotter och barnbarn har bilproblem, och den stackars lilla flickan ser varm ut i hettan.
En kvinna kittlar en man på golvet medan fem andra skrattar.
Tre herrar som använder en slang för att pipa ut något ur en oljetrumma.
En man ger två tummar upp till en massa människor.
En slaktare skär kött i en affär på disken.
Man och kvinna dansar en solig dag på en gata kantad av små byggnader och utomhusutställningar.
Ett plan flyger ovanför medan en man går nära vattnet på en strand.
Unga vuxna dansar på gatan
En flicka i en ljusgul jacka står framför en ljusgul lastbil.
En vaktmästare sopar trottoaren på en livlig gata med många bilar och fotgängare.
Två unga bröder, klädda i uniform, övar kampsport på föräldrarnas balkong.
Några personer sitter tillsammans på den snöiga bergstoppen.
Två män sopar ett rum som är tomt förutom en stege.
En man sitter i sitt tält på ett berg.
En svart hund är redo att fånga en frisbee.
Barn fördriver tiden medan andra tittar.
En man står i en röd skjorta och blå jeans mot en man i svart över spåren med en rulltrappa i bakgrunden.
En man och en kvinna dansar medan åskådare tittar.
Ett band spelar utomhus spelar gitarrer och trummor, sångaren bär solglasögon och en svart skjorta och bandanna med en getmö, den andra mannen bär en fedora och lila skjorta, de andra spelarna är inte avbildade.
En ung musiker uppträder framför en skyline.
En arbetare med randig skjorta och handskar som håller fast hans hatt med ena handen och skrevet med den andra.
En man i formell klädsel spelar klarinett
Två män rider cykelspår och hoppar över en kulle i ett skogsområde.
En ung man i blå skjorta är i luften med en cykel
En bicyklist som bär en ljusblå kortärmad t-shirt och skyddande ansiktsväxel utför ett trick där han är helt upp och ner, inramad mot en bakgrund av barrträd och en delvis molnig himmel.
En man som grillar utomhus med några personer som njuter av hans kött.
Vissa män och pojkar leker med en frisbee i ett gräsigt område.
En man poserar ser tillbaka medan en yngre flicka fiskar.
Ett asiskt barn med en gul rosett i håret på en sving med en asiatisk kvinna som står bakom henne.
En liten pojke med en fotboll som flyger.
En ung dam på ett gymnastiskt evenemang mitt i sin föreställning, klädd i en blå och vit dräkt medan lagkamrater tittar på.
En man övar med en tredelad stab framför en röd gardin.
En man klädd i en ljusblå skjorta dumpar saker från en soptunna till en annan soptunna, medan han står i ett rum fullt av matdonationer.
Barnen går längs en grusväg.
Två postarbetare ler medan de håller soptunnor med konserver.
Ett litet barn som leker i en Lexmark box och använder den som ett fort.
En balettdansare i en blå leotard som gör en ryggböj med sin vänstra hand utsträckt.
En liten pojke i orange skjorta med flip-flops har handen på huvudet.
En man i grå skjorta som spelar visselpipa.
En sjuksköterska lyssnar på en annan kvinnas hjärtslag med ett stetoskop.
En kvinna med brunt hår gör ett vetenskapligt experiment medan hon bär glasögon och en blå skjorta.
En liten unge i blå rock som tittar på ankor som simmar.
En man i våtdräkt surfar på en vit surfbräda.
Hunden hoppar i snön nära ett träd.
Fyra pojkar visas i ett hus som leker och alla bär t-shirts.
Två män i hårda hattar sågade en planka av trä.
Tre män sitter på en båt och tittar upp mot himlen.
En nunna ger en man en servett.
Fyra dansare klädda i vita, flödande klänningar utför sina rutiner.
En ballerina i röd klänning hoppar upp i luften.
En kvinna ger dockor från ett stort fönster till en annan kvinna utanför på en stege.
Det finns fyra soldater, två skadade och i rullstolar.
En man som spelar på en basebollmatch som just har slagit slagträt.
Folk som står utanför och väntar på att graffititåget ska passera.
Tre kvinnor klär ut sig till ninjor för en maskerad.
Ett barn i en vit skjorta som klappar händerna.
En man i röd tröja och blå mössa målar en bild.
En kines spelar trummor i ett band.
En asiatisk kock som bär vitt skär kött på en restaurang.
Män i köket lagar mat.
En liten flicka i blått tittar på en liten pojke i svart sving på en disney prinsessa pinata.
En liten flicka med ansiktsmålning som svänger en pinne på en pinata.
En äldre man som bär en solbränd tröja arbetar på en målning.
En gammal man i röd jacka håller upp pengar.
En kaukasisk kvinna hoppar och slår ihop sina klackar inför en skara afrikanska barn.
En man och en liten pojke njuter av en middag med grönsaker.
En tonåring fyller sin mun med något när han sitter inne i ett hem.
En man spelar dragspel.
En man med halsduk kastar en stickspätta på en övergiven strand.
En man i hatt och blazer uppträder på gatan med sin gitarr och munspel.
Två män böjer sig över de hydrauliska slangarna på en John Deere-anläggning.
Två kvinnliga gatuartister interagerar lekfullt med en boll som rekvisita.
En amish dam hänger upp kläder för att torka ute på en linje.
Två unga flickor visar fingeravtryck på en linjeteckning av ett djur.
Den lille pojken vadar genom poolen med röda armfloaties.
Det finns en grupp människor som spelar fotboll bredvid ett gäng cyklar.
En man i vit hård hatt drar en havssond som lyfts över båtens sida.
Två små pojkar rode sig genom det bruna skumma vattnet.
En liten pojke hoppar högt ovanför poolen med en man i bakgrunden.
En pojke bär baseballhandske och håller i en baseball.
En grupp människor sitter på en bänk och beundrar en målning i en utställning medan andra går förbi.
Crowd rör sig genom byggnaden med stora skulpturer centrerade i bild.
En man med ryggsäck, bär shorts och en t-shirt, går genom ett konstmuseum, tittar uppåt.
En man och fyra tonårspojkar räfsar en baseballdiamant.
Studenten använder en kamera för att ta en bild av ett konstverk.
Eleverna är noga fokuserade i en riktning.
Inomhus fungerar en kvinna som bär kirurgisk mask, klänning och handskar på en person som lutar sig tillbaka.
En grupp killar som jobbar som grupp i ett klassrum.
En man skateboards i en skatepark medan andra åkare skakar i bakgrunden.
En man och ett litet barn leker ute i gräset.
En lastbil med en kran och 3 anställda på den är framför ett byggprojekt som har en grön beläggning.
Ett litet barn kastar en frisbee till marken.
Indiska kvinnor lär sig av en man hur man tillverkar tyg.
En man är klädd som en filmperson som håller en pistol i lobbyn på en biograf.
En polis sätter koppel på en hund.
En polisman rider en häst genom gatan.
Många kvinnor försöker och tittar på bärbara datorer i en Walmart.
En manlig tennisspelare förbereder en vänsterhänt förhand medan han spelar på lera.
Den gröna hulahoopen svävar genom luften när den unga damen tittar på när den landar.
Mannen i rött står bakom kedjorna medan han tittar över vattnet mot land.
Nio män spelar kraftfullt rugby på en utomhusplan.
Två män slåss inför en folkmassa.
Odd barn med falska ögon barrows och ett snitt på läppen håller ut sin högra hand.
En kille som sitter utanför på en hink och spelar banjo.
En tennisspelare gör sig redo att slå bollen medan man står på en ljus orange bana.
Två honor klädda i rosa sitter på gungor som är en del av en upphängd trä fyrkantig vara.
Två barn tittar genom ett teleskop på en gata i staden, och pojken använder en stegstege för att se igenom glasögonen.
En grupp barn i vattnet håller upp en blond pojke i röda badbyxor.
En man visar några lådor med parfym för en person inuti en bil.
Barn leker utanför.
Två kvinnliga armépersonal hanterar mycket pappersarbete vid ett skrivbord.
En kvinna gör hantelpressar på ett gym.
En kvinna i en svart och vit rutig skjorta färglägger i en färgbok med en liten blond tjej.
Grupp av människor vid havet som innehar ett nät
En grupp män och kvinnor sitter vid ett restaurangbord med öl och mat.
En ung kvinnlig baseballspelare glider till hemmabas men fångas av umpiren.
Två personer hoppar på en bro i bergen.
Kvinnan, i den blå skjortan, bär en kvast och en metallstoft.
En liten flicka går vid stranden i blå och röda regnstövlar.
En blond liten flicka tittar genom en grön kikare.
En pojke klappar en hund på en gård med en trädgård i.
Brunhåriga kvinnor presenterar födelsedagstårta för blondhårig pojke framför publiken.
En grupp människor i alla åldrar samlas i ett ganska vitt kök för förfriskningar.
En ung pojke och en kvinna poserar nära en snögubbe som en hund ligger på den platta, snötäckta marken.
En liten pojke i flanellpyjamabyxor och en orange skjorta spelar gitarr på soffan.
En pojke är täckt av sand på stranden.
Ett barn bär grå byxor, grön vinterrock och svart skidmössa matar gäss i en sjö.
En man målar en vägg.
En ung pojke kör sin pedaldrivna leksakstraktor utomhus när hans vän hoppar runt i bakgrunden.
Ett barn i en röd snödräkt står bredvid en snöhög.
En pojke och flicka står tillsammans, och flickan håller i en volleyboll.
En liten flicka och pojke leker te med låtsasrätter och dockor vid ett litet bord.
Två små barn klädda i vinterkläder rider sina leksaksslädar nerför en liten kulle.
En byggnadsarbetare i orange väst sträcker sig över arbetet.
En kvinna och en manlig barn är engagerade i en ballong kamp som en man tittar på.
En tjej i blå klänning leker med en kinesisk jojo.
Tre unga kvinnor i vita och svarta klänningar spelar fioler på en scen.
Ett barn använder en hand för att radera en del av en annons från en krittavla.
Två personer, en med blå skjorta och en med rosa skjorta, rycker ner en byggnad.
Två arbetare som jobbar på ett tak och tittar över en stad.
En man håller en kvinna i en blå och vit dräkt i luften.
En militär grupp marscherar framför en McDonald's
En entusiastisk liten flicka som visar sina färdigheter på trummorna.
En spelare på stranden väntar på att fånga en boll.
En manlig fotograf knäböjer medan han tar en bild med en Nikon kamera på en parkeringsplats.
Två kvinnor har en diskussion på ett mestadels vitt, modernistiskt kontor.
En stor skara människor, och vid sidan av en gentleman att få sin bild tagen av en fotograf som han poserar.
En affischtavla för Comcast Digital Voice som refererar till Madagaskar 2.
Ett barn i röda och blå floaties tittar ner på vattnet.
En äldre man som plöjer en gitarr i ett band.
En kvinna håller två små flickor medan hon sitter korsbent på gräset.
En hjälmhjälmad bergsbestigare stiger upp på en klippa med träd bakom sig.
Flera små flickor klädda i kostym för att underhålla sina vänner och familjer.
En flicka hoppar rep på en parkeringsplats.
En grupp människor står i kö utanför Hyatt Regency.
En tjej med blå höjdpunkter ser en hund hoppa för att fånga en frisbee.
En liten flicka hoppar rep på en parkeringsplats.
En kvinna spelar ett tangentbord medan hon sjunger in i en mikrofon.
Två byggnadsarbetare manövrerar en stock på eller av en plattbädd på en kraftigt trädfodrad väg.
En man i hängslen dansar på en scen medan ett band spelar bakom honom.
En man står på en bergstopp och tittar i fjärran.
Barn leker på trottoaren omgiven av löv.
En manlig vandrare bär sin utrustning uppför det snöiga berget.
En man som åker skidor i bergen
En man står på toppen av ett berg och stirrar på solnedgången.
Ett barn observerar ett exemplar i ett mikroskop.
En ung flicka i svart går på ett löpband.
En grupp människor som tränar på ett grönt fält.
Män och kvinnor utövar yoga i en offentlig park.
Två kvinnor med kjolar dansar på en scen.
En man som pekar mot publikområdet på scenen medan han håller en mikrofon med banjos bakom sig.
Två kvinnor möter varandra i en dans.
En grupp rullskridskor följer en man som bär blå byxor och en röd skjorta på ett träpanelgolv.
Två bruna hundar leker med en röd boll.
En ung man i en baklänges basebollmössa balanserar sin skateboard på kanten av betongen.
Den unga damen står upp efter att ha spelat i en pjäs.
En kitesurfare och en drakflygare förbereder sig för att lansera sina respektive drakar på en gräsbevuxen sluttning.
Barn som leker på en lekplats med en man som sitter på en bänk och läser en tidning.
Två kvinnor går på en grå väg.
En man i kostym och hatt håller ett vinglas.
En baseman håller ut sin handske för att fånga en boll och tagga ut motståndaren.
En kameraman jobbar på ett sportevenemang.
En kvinna i en turkos topp som pratar med konduktören av en vagn nära ett utländskt café.
En man i en blå skjorta tvättar ett fönster högt från marken.
En kvinna med grönt hår, en sexig outfit och svarta stilettostövlar står i en pos bakom några svarta räcken.
Tre människor rider hästar är i ett lopp.
En stor skara människor höjer sina armar i en urban miljö medan fotografer dokumenterar händelsen.
Ett litet barn som dansar framför ett orkesterband.
Män och kvinnor som äter nära en butiksyta en man och en kvinna med en barnvagn som tar till varandra.
Ett barn med blont hår stirrar in i en kamerabild.
En ung kvinna med en fjäder i håret finns bland en skara människor.
En cowboy på en häst på en rodeo.
Asiatiska religiösa medlemmar bär mörkröda kläder är på en utomhusmarknad samtalar med beskyddare av en grönsaksstånd.
En liten pojke som hoppar i en stor vattensamling.
En simmare simmar från ena sidan av poolen till den andra.
Fyra män sitter på en bänk i en ökenby.
En kvinna i gult arbetar på ett fruktstånd utomhus medan en kund i solglasögon står nära montern.
Grafik Designer, manlig (ungefär 38 år gammal) utformning på designbordet på kontoret.
En man i svart och vit dräkt och bär en svart hatt och vita handskar sitter på en förstärkare och spelar en tuba med lågor som kommer ut ur öppningen.
Unga dam under en föreställning av modern dans.
Ett barn i grön skjorta tittar på något som är utanför ramen.
En flicka, i en rosa skjorta, njuter av en utsökt godbit sockervadd.
En kvinna i en flytande grön klänning dansar.
En gentlemän njuter av en eftermiddags golf.
En svartklädd man spelar ett långt instrument med andra i en orkester.
Tre kvinnor i träningsoveraller, böjda över, städa en basketplan.
En man klädd i rött och gult rider en röd sportcykel kör på en kapplöpningsbana.
En man sitter på en pall och läser en tidning på en trottoar.
En krulhårig hund försöker bita en annan hund i en grön och orange krage.
En stor grupp människor står i två ovala medan de lyssnar på ett bandspel i bakgrunden.
En kvinna i dykutrustning skrattar när hon står nackdjupt i en simbassäng.
Folk tränar i en studio med kuddar.
En kvinnlig sångare på scen med en tamburin med två män som spelar gitarr och trummor.
Rodeo ryttare visar bra stil mitt i hopp av hans bucking häst
Två kvinnliga tennisspelare skakar hand över nätet medan en tjänsteman och hovvakt tittar på.
En cowboy rider en vild häst men håller knappt fast vid en rodeo.
En flicka klädd i svart hoppar i luften medan hon håller i snöret på en rosa ballong.
En liten flicka som springer genom en massa människor som sitter.
En brudgum klädd i en svart smoking doppar och kysser sin brud vid bröllopsmottagningen i ett hem.
Flera människor dansar i ett trångt rum.
Mannen i en blå skjorta med ID-brickan dammsuger en modell av en byggnad.
En orientalisk man i vit skjorta som säljer mat utanför.
En man sitter ovanpå en gatubelysningsstolpe med en bild av en sak i ben som ser upp till honom i fokus.
En grupp män, en med cykel, på en brygga med däck och rep.
Två män arbetar i ett fält av en håla som deras hund är på väg att gå upp på dem.
En pojke utför ett stunt på en skateboard i en skatepark.
En grupp män står runt ett bord och tittar på en karta.
Baby har kul att borsta tänderna.
En kanna i en blå skjorta, på högen, övar sitt grepp innan han kastar planen.
Baseballspelaren är på väg att springa på en bas.
En basebollspelare svänger på planen medan motståndarlagets catcher är redo för bollen.
En man i en vit baseballuniform som plockar upp en baseball.
En bas löpare är taggad ut av motståndarlaget.
En man i baseballkläder försöker fånga baseballen.
En baseballspelare i en röd och vit uniform ser på som hans lagkamrat resor medan du springer till en bas.
Spelare 22 får tonhöjd från kvinnor nära kannor mount.
En man i en rutig rock säljer färgglada ballonger från en vagn när folk går förbi.
Ett barn tittar ut genom fönstret på en buss.
En liten pojke i grön skjorta leker i vatten med en liten flicka i rosa skjorta och lila kjol.
Människor går och står runt en stor fontän, två barn står framför fontänen.
Tre killar på scenen, varav en har en gitarr och en annan ett tangentbord.
Två pojkar leker i sanden.
En äldre kvinna som bär förkläde och svart klänning hänger kläder på tvättlinan.
Unge pojke spelar ett spel på datorn.
En man i en gul tanktopp kör en traktor med flera passagerare.
Skolbarn i uniform sitter på kullen, medan de äter lunch.
En konditorikock strör ingredienser på en kastrull med bakverk.
Några barn och vuxna som har förkläden på sig och bakar kakor.
En man med en galen frisyr och en lång flätad mustasch sitter på trottoaren utanför och spelar ett stränginstrument.
En kvinna och en flicka tittar på en svävande boll tillsammans.
En liten pojke i blå mössa och blå skjorta tittar på en modell medan han står utanför.
Man skär upp sin mat för att sätta på en tallrik.
En grupp multietniska ungdomar sitter i en cirkel på gräs bredvid en kulle.
Ett par som håller varandra i handen när de går nerför stranden.
Ett nygift par poserar för formella bilder framför en vacker vattenfontän.
Ett hejarklacksteam av unga flickor uppträder på en utomhusplats.
Sex män i gula kostymer och orangea livvästar lämnar en stenig strandlinje på sin båt.
En person sitter i stenar i vattentät utrustning med sina stövlar i vattnet.
Tre personer försöker känna ruset av fritt fall innan de drar sina fallskärmar.
En ung pojke tittar på en man målad i allt guld.
Mina herrar som sitter i en halvcirkel och spelar mässingsinstrument i parken
Män i Amerikanska Revolutionära hattar och kostymer står med amerikanska flaggor, baklänges till kameran.
En tjej och en kille som ser ut som de är utanför breakdancing.
En man som bär på en blå oljetrumma utför en show på gatan.
En man bär amerikanska flagga shorts, skjorta och hatt vid en utomhus sammankomst.
En man är på väg att träffa vattnet.
En grupp människor samtalar medan en man i vit skjorta antecknar.
En grupp män håller ett möte.
Kannan på högen, nummer 46, är redo för nästa pitch.
En basebollspelare, klädd i rött, dyker för att fånga en boll.
En basebollspelare i blått märker en spelare i rött ut.
En kvinna med grönt hår hula hovar inför en folkmassa.
En ung flicka med blont hår som kikar genom ett mikroskop.
Kvinnor i svart rock väntar på tvätt medan de läser tidningen.
En man sitter i sin stol på ett kontor medan han sätter på sig en röd fleecetröja
En äldre man spelar gitarr medan han är på scen.
En man och en kvinna skapar en matsal.
En man deltar i en uråldrig rituell dans.
En man i blå jersey och röd hatt ska kasta en baseball.
Tre män jobbar på en byggarbetsplats.
En baseballspelare som glider in i hemmet som motståndarlagets catcher väntar på baseball för ut.
En baseballspelare med en röd hjälm träffar en baseball.
Afrikansk livsmedelsmarknad, med dam shopping för grönsaker och frukter.
En ung flicka blåser en stor bubbla på sin veranda.
Flera män i vit kockjackor arbetar i ett kök.
En tjur springer mot en röd duk.
En död tjur dras ut från en arena av hästar.
En person med långt hår sitter på en lila soffa.
En man med ryggsäck på väntar på vid en deli disk av en kontorist med svart hatt.
En grupp människor går uppför en sluttande stig kantad av träd.
Åtta unga kvinnor utför en hejarklacksdans på en domstol.
Mannen i den vita skjortan ber offentligt.
Person i vit skjorta och blå jeans, håller handen ut med en tom kopp i den andra, och en flytande röra på marken.
Långa köer väntar på att få komma in på The Magpie Cafe.
En skjortlös man är i luften med en skateboard under sig.
Individer sitter förnöjt på parkbänkar under nyblommiga träd i ett urbant område.
Två kvinnor är på bankomater och får pengar och damen till vänster har två barn.
En man tar bilder på sin telefon av stenfigurer medan hans hund tittar på.
Ett ungt par som rider på en buss med pojkens arm runt flickan.
En liten pojke går genom skogen.
Folk rider en rulltrappa upp och ner för en tunnelbanetunnel.
En kvinna uppträder en infödd dans framför ett band.
En kvinna i etnisk klädsel knäböjer på marken och böjer ryggen i en dansposition.
Fyra personer har svarta leotards som dansar på en strand.
Tre barn på nära håll på stranden med fler människor i bakgrunden.
Folk njuter av en trevlig omgång bowling.
En mystisk man lutar sig mot den vita väggen i en svagt upplyst tunnel.
En man är på en tjur på Rodeo.
En svart kvinna kikar genom ett teleskop med flera personer i bakgrunden i parken.
En man tittar på månen kastar ett teleskop i skymningen.
Två asiatiska män sätter sig ner och tittar på något som inte syns på fotografiet.
En ung överviktig hane ställer upp en boll.
En äldre vit man med glasögon arbetar med ett metallarbete på ett städ.
Tre byggnadsarbetare som fullbordar grunden för en uppfart.
En dam som bär röd hatt fiskar i en lugn och fridfull sjö.
En kvinna i klänning hängande tvätt uppe på en klädstreck utanför på hennes gård.
En ung kvinna målar väggen i ett rum med klar orange-röd färg.
En man pressar någon sorts degliknande mat mellan två träpaddlar.
En kvinna, med mörkt hår i fläta, som ler som en grupp duvor flyger runt henne.
En man kör förbi en lastbil som kör fordon.
En man med grå skjorta med taggen bombardier använder en orange ficklampa.
En grupp arbetar med ett pianoprojekt och har 53:11 kvar.
En grupp människor med vitt ansikte smink samlades runt ett bord med vissa människor spelar instrument framför en lastbil i bakgrunden.
Det finns en snickare som mäter ett bräde.
En man i grå tröja och glasögon skrattar.
Kontortionist i underlig rutig outfit klädd i vit mask.
En brunhårig kvinna ger en svart och vit hund en frisyr.
Man bär en hård hatt och ansiktsmask medan man står sysslolös på jobbet.
En man längst ner i ett betonghål med ett rep.
Två kvinnor som bär skyddsglasögon, tittar på samma anteckningsbok.
Män samtalar som två män är i en hink hiss.
Kvinnor njuter av en dag shopping på gatorna.
Kvinnor dansar i ljusa kostymer och bara fötter.
En fågel syn på kvinnor som dansar med olika färgade klänningar.
Fyra tjejer synkroniserar dansscener där de bär blå och lila kläder.
En liten liga kanna kastar bollen
En kille försöker göra en bas och den andra kastar en boll.
En sångare knäböjer med sin mikrofon medan en trummis spelar i bakgrunden.
En man som lutar sig över ett stängsel pratar med en baseballspelare som vilar.
Pojke hoppar från den höga dykarbrädet vid en allmän pool.
En jockey hukar lågt och driver hästen framåt under en hästkapplöpning med en annan jockey i het jakt.
En häst jockey täckt av lera under ett lopp.
En jockey på en vit kamel tar ledningen i en kamelkapplöpning.
Tre unga, atletiska flickor är klädda i svarta och blå leotards.
En kille med blå jeans på och några i bakgrunden städar upp en stor röra.
En massa människor som ser en man cykla på en smutscykel.
En man i blå påfågeldräkt med rök och dimma under sig.
En basebollspelare som fångar en boll när det kommer till honom.
En tjej i slitna jeans och en vit t-shirt leder andra i en synkroniserad dans.
En asiatisk gymnast i en Rheinstonedräkt som håller i en batong.
En manlig skateboardåkare i svart skjorta och vita byxor som hoppar över ett gult föremål.
Fyra unga flickor tävlar i laggymnastik.
En ung gymnast i en bourgogne och silverleotard utför en rutin.
Det finns en kille som gör tricks med sin skateboard.
En kvinnlig gymnast gör en flip som fångas på fotot med fötterna i himlen och han går mot marken.
En man använder ett paraply.
Två pojkar sköts av en vattenpistol av en annan pojke på en gård.
Indianerna har en samling med rockar och mat och dryck.
Under en vattenstrid bestämmer sig en pojke för att fördumma en liter vatten på en flickas ansikte.
Ett band framför musik på en scen med ljus.
Blond man i svart kostym med gula skor i hoppning över ett hinder.
En åsna upphängd i luften efter en vagn den är fäst vid över varv.
Två män slåss mot varandra i en kampsport match.
En person i en orange kajak navigerar vita vatten forsar.
Två män kör motorcykel med ett fack på sidan
En fullsatt torg som underhålls av gatuartister.
Två män arbetar på flickor cykel framför garaget.
En medelålders man i röd kostym fixar sin cykel.
Två marinsoldater och två unga flickor har monopol.
En man står i en tvättstuga och pekar på en knapp på en tvättmaskin.
Två pojkar i ett skogsområde placerar löv i en klar utsiktsbehållare.
Två musiker uppträder på scenen inför en publik.
En man i skinnjacka som håller en hjälm på en trottoar.
En man gör en kanonkula i en pool, stadion stolar fyller bakgrunden.
En kvinna klädd i neonrosa tutu och leotard håller dramatiskt sina boxningshandskar ovanför huvudet i ett trångt offentligt rum.
Fem personer står på en modern rockkonsertrepetition.
En liten pojke håller en basketboll i position att kasta den i en båge på ett spel.
Tre simmar konkurrenter med blå, gröna och gula huvudmössor gör sig redo att tävla.
En tonåring i en blå t-shirt i att spela ett spel vid ett bord vid en video arkad.
En man som spelar synthesizer med grön tröja och hatt.
En fotograf i grön skjorta och jeans, stops för att fotografera en simmare i rött som lämnar poolen.
En kvinnlig idrottsman springer efter att ha lämnat en simbassäng.
En ung flicka äter en tårtbit.
Män tävlar i en motorcykeltävling.
En skjortlös man i svarta byxor drar benet på en annan man i gröna byxor.
En baseballspelare hoppar mot stängslet för att göra en fångst
En baseballspelare i vit uniform kastar bollen till en annan spelare vid en bas.
Två män spelar cricket i en park.
En baseballspelare i grå uniform fångar en boll i sin handske.
En pojke spelar på en grön gunga.
Ett gäng glada barn som har kul badar och en pojke visar upp sin talang med en back flip.
En kvinna med rött hår sjunger.
En flicka i rött med en vit tutu utför ett danssteg medan 6 andra flickor står bredvid henne.
En trött man i en blå skjorta paddlar nerför en sjö.
En man med hatt på vid havet, lyfter upp en säck.
En person i rosa försök att montera en häst.
På en rodeo, en brash cowboy har vred en ung kalv med många fans i bakgrunden tittar på dem
Simningskonkurrenterna förbereder sig för sitt möte.
En baseballspelare i vitt glider in i basen medan spelaren i grått försöker märka honom.
En motorcyklist som utför fantastiska trick framför tusentals människor.
Två hundar leker tillsammans på gräset framför en liten stenbrunn.
Anställda försöker fixa de trassliga näten till fiskebåten.
Två män sitter på en hög med fiskenät på en brygga bredvid ett noggrant utformat fiskefartyg.
Ett band spelar för en krona i en nattlig miljö.
En man som bär en grön skjorta spelar musik på en blå uppsättning trummor.
En åkare som rör sig runt ett spår framför en publik.
En man på en skatepark gör en Ollie ur en skål nära en strand.
En tjej klättrar över en massa kablar.
Baksidan av två män som lagar mat vid en spis.
En man vänder sig genom luften med en stor tall i bakgrunden.
En pojke dansar med hörlurar i örat.
En man i vit skjorta som blåser i trumpet.
Kvinnan försöker surfa framför två fotografer som tar bilder.
Den här kvinnan rider på en solig eftermiddag.
En person som rider på en gruscykel farligt nära en klippa i en skog.
En man och en kvinna på hästryggen som håller upp den amerikanska flaggan inför en rodeo.
En ung pojke i en blå t-shirt tittar genom ett mikroskop.
Två kvinnor deltar i antingen beredning eller försäljning av något i gula påsar.
Tre män spelar musik på en scen, en är på pianot, en sjunger, medan den andra spelar en trumma med händerna.
En surfare som visar upp sin talang offentligt med hjälp av en konstgjord vattenmaskin.
En kvinna läser en tidning när hennes tvätt blir klar.
Fyra nakna pojkar leker med en oxe i smutsigt vatten.
Det här är en man i clownkostym som balanserar ett tefat ovanpå en pinne, på näsan.
Tonåringar som spelar gitarr live i ett rockband
En dam tittar på en blå låda medan den kortare damen tittar på något på sin telefon i mataffären.
En roller derby matcha med en actionbild av en derby flicka i förgrunden.
Två damer i tank toppar sjunger in i en mikrofon, de båda har mörkt hår och den ena är vit och den andra afroamerikanen.
Två dykare inspekterar ett stort metallföremål i vattnet.
En man som spelar gitarr på scenen under rött ljus.
Flera honor sitter indisk stil gör vad som verkar vara textila arbete.
En kvinna i blå skjorta talar med två andra kvinnor och en man, som bär glasögon.
Två män jobbar med dator-DJ-utrustning i mörkret.
En kvinna kör ett hjulförsett föremål med en ponny på framsidan vid en strandpromenad.
En grupp barn och unga vuxna som åker skateboard på en ramp.
En grupp av turister på en liten båt med byggnad runt som är omgiven av vatten.
Ett par sitter tillsammans vid ett litet cirkulärt bord i en äldre, rustik byggnad.
Två båtar med paddlare och passagerare är i en flod kantad av byggnader.
En man som ger en presentation medan han bär en brun randig kostym.
En man som bär solglasögon och hatt står på ett fält av vilda blommor och inspekterar en av blommorna.
En upptäcktsresande på en grusstig som tittar på en blomma.
En person som bär en mössa och en blå rock står böjd över resväskor av olika föremål, inklusive kameror och saxar, på trottoaren.
Flera män på däck på ett skepp sänker ner en annan man i vattnet.
En man som sitter på golvet ser ut genom ett stort fönster.
En man gör ett enhänt handstöd på ett trägolv.
En man får ett papper från en kvinna medan hon skakar hand, när en man som bär en "Ohio State Geografi" skjorta ser på.
Två män i karateutrustning med stridspinnar.
Mannen är ivrigt håller upp en fläktad kortlek av spelkort.
Någon viskar ägg med en handhållen mixer.
En man använder sprayfärg för att måla en bild på en vägg.
En man balanserar i en pose som en kvinna springer nerför kajen vid honom
En kille med svarta kläder gör balett framför piren där man kan se ett kryssningsfartyg.
Mannen i svart poserar för en bild.
En man klädd i svart på stranden som sitter under ett rött paraply.
Familj och vänner väntar i närheten medan en grupp tar en simtur vid inomhuspoolen.
Den här mannen verkar omedveten om insekterna som liftar med honom och hans vapen.
En man klädd i grått liggande på golvet framför en annan person medan han sträckte ut handen.
En person flyger genom luften fäst vid en bräda med en fallskärm.
Det är en kvinna som borstar tänderna i skogen.
En cyklist som gör ett trick från en ramp som lyder "RONA" och "Cariboos Brewing".
Folk är i en tvättmatta och tvättar kläder.
En man som bär heta rosa kalsonger står på en utomhusplattform och jonglerar framför en publik nedanför.
En man som bär hjälm och kör en fyrhjuling som visar upp sig för kameran.
Flera åskådare tittar på när en man gör en wheelie på en gul fyrhjuling cykel
En ung man sparkar en annan ung man framför ett tvåvåningshus.
Denna vackra dansare sträcker sig i en studio, antingen värms upp eller kyls ner.
En kvinna med ett målat ansikte håller en fläkt framför ansiktet.
Ett barn ser ganska trött ut när hon sitter inne i en bagageväska.
En kvinnlig kock visar upp sina snidade frukter.
Gubben skär en bit rör till rätt form.
En matsalsbil för skådespelare på plats som filmar ett stycke om 1800-talet.
En arbetare i orange väst och hård hatt är ovanpå en gul stege som arbetar på en telefonlinje, medan andra män arbetar under.
En snåljåpare utför ett trick i vattnet.
En person står i en båt märkt Texas Mooring framför en röd vägg.
Framför en klädaffär lägger en man tegelstenar.
Ett litet barn sätter sig fast i en sten på stranden av en damm med en hund i närheten.
En ung blond pojke leker med ett dockhus.
En kvinna sitter vid ett skrivbord och skapar halsband av diverse pärlor för hand.
Isuzu lastbil kör förbi medan en man med några kor kör motsatt väg.
Ett litet barn cyklar bort från en stor bro en molnig dag.
En grupp män sitter längs en blå vägg bredvid två cyklar som bär korgar med frukt.
Tre barn leker med en volleyboll i grunt vatten medan en vuxen i en röd mössa och neongrön skjorta observerar.
En tatuerad man i en tanktopp skriker in i en mikrofon.
En man och en kvinna på cyklar cyklar nerför en stor motorväg i leden körfält, tillsammans med andra cyklister och joggare.
En liten pojke tittar på några föremål genom ett förstoringsglas.
En kvinna i orange skjorta hänger kläder på en klädstreck utanför.
Ett barn står i högt gräs vid en vattensamling.
Dam i grå topp och vita byxor bär tvål i tvättmatta.
Hunden på bilden gillar inte att blåsa torktumlare.
Två män bär traditionella skotska kläder, håller säckpipor i sina händer.
En man jonglerar med flaskor som brinner.
En tennisspelare, bär en gul skjorta, hoppar för att träffa bollen till den andra spelaren, som bär svart.
En ballerina dansar i en mörk, rustik miljö.
En skjortlös man är bergsklättring i en mycket brant vinkel.
En kvinna som står bakom en flicka och hjälper flickan med ett experiment.
Två kvinnor i vita skjortor står vid ett handfat, en med en skål och en med en penna.
Forskare ser vätska flöda ur en bägare i ett labb.
En man i en labbrock gör något slags experiment i ett labb.
Två joggare och två cyklister vill ha plats på den här gatan.
En kassörska som står framför kassan med pengar i handen.
En man i en lysande grön skjorta står på en trottoar.
En mycket ung pojke sitter på sin förskolecykel under ett utomhusbord.
En man i flottan letar efter nåt.
En ung flicka med mörkt hår böjer sig över ett lerkärl som ligger på ett bord.
Det finns en flicka som skapar konst i den här bilden.
Folk beställer fisk på vad som ser ut att vara en asiatisk fisk- och skaldjursmarknad.
En ung man i randig skjorta med gasmask på.
En arbetare använder en hammare och mejsel för att göra sniderier i trä.
En man arbetar på en restaurang medan en man diskar bakom sig.
En skallig man i vit skjorta knäböjer på en träplattform och tvättar huvudet i en bäck.
En grupp människor, allt från barn till vuxna, som förbereder sin utrustning innan de dyker.
En man i hatt lutar sig mot en delvis byggd träkonstruktion.
Ett harmoniserat ögonblick i en färgglad ballerinashow.
En grupp rullskridskor åker skridskor på en bit cement med palmer i bakgrunden.
En pojke med hjälm mountainbikes genom skogen.
En kvinna som spelar fiol med solglasögon på huvudet.
En man räddar en annan man från en båt.
Två män i polisuniform pratar.
Tre personer, två män och en kvinna som spelar domino på ett runt träbord.
Asiater dansar på gatan med träd och byggnader i bakgrunden, medan de bär röda, vita och gröna dräkter med gröna pannband.
En grupp asiatiska människor i dekorativa klänning leende, och gå lyckligt i en parad.
En laboratorietekniker undersöker ett blodprov med hjälp av ett högeffektivt mikroskop.
En gammal man och unga kvinnor som dansar på en fest.
Två poliser sitter på motorcyklar på vägen.
En blond kvinna spelar gitarr på scenen.
En cowboy försöker att inte ramla av den böljande ko, medan åskådare, en man på en häst, och en rodeo hjälpare observera.
Tjuren spottar när männen försöker lasso den.
En man skär träplankor med en bordssåg medan en annan man tittar.
En man i orange uniform står mitt på gatan.
Bandmedlemmar marscherar i en parad på en trädkantad gata.
Tre vandrare går uppför en brant kulle i ett vackert skogsområde.
Folk balanserar på bjälkar som kommer ut från en John. F Hunt ägde Genpac generator.
En grupp människor vandrar längs ett gräsområde.
Två unga flickor sitter på en trottoar färg på det med krita
Två personer står i havet och håller ett nät medan den tredje personen tittar
En musiker på gatorna bär shorts och stylar en mohawk.
Fyra personer ro i en kanot på en lugn och fridfull sjö.
En grupp unga människor som bär baddräkter står på en klippa över vattnet, och en av dem är redo att hoppa i vattnet nedanför.
En liten flicka och en kvinna som borstar tänderna.
En mor och två små barn sitter på en soffa utanför trottoarkanten.
En man på en mobiltelefon får sina skor lysta av en annan man i blå uniform.
En långhårig, skjortlös man med ansiktsfärg spelar en basgitarr på en konsert.
Ett djur försöker korsa floden.
En man i grön skjorta bär en flagga mitt ibland en grupp människor.
Arenan är fylld med åskådare som tittar på ett sportevenemang.
Många människor på ett byte träffas på en parkeringsplats.
En fotbollsmatch spelas.
En kvinna bowlar barfota som 2 personer i bakgrunden huvudet mot videospel.
En liten flicka ligger på en matta, färgläggning.
En publik som bär orange hejar på sitt lag på en stadion.
Fem personer går över ett idrottsområde, en man bär älghatt.
En man bär en blå och gul racing uniform samtidigt hålla en flaska
Ung pojke möter andra barn, också rider cyklar.
Ett spel av Carcassonne spelas på ett bord medan en kille överväger sitt drag.
Den unga flickan leker glatt i trädet.
Två pojkar, en i vitt och den andra i brun skjorta, spelar ett tv-spel medan en tredje tittar på en väska.
En man i svart skjorta som äter god mat.
Ett inbördeskrig med kanonteam som avfyrar kanoner.
En kvinna som bär huvudduk arbetar med sina händer.
En pojke i en skatepark som bär en blå hjälm inline skridskor på ett litet räcke.
Ett fotbollslag spelar, det gula laget har bollen.
Två män, en klädd i officiella kläder, står på en båt.
Mycket fattiga människor i ett främmande land spelar ett spel för att underhålla sig med vad de har.
En publik samlas och hejar på en scenföreställning.
En ung kvinna som bär cykelklädsel vänder sig bakåt
En kvinna med tennisracket böjer sig ner, med graffiti i bakgrunden.
Ett barn som bär en piratdräkt håller upp en skalle och korsbensskylt.
En tjej i blå skjorta sitter i en salongstol och får håret gjort av stylisten.
Barn i röd skjorta väntar i linje med många andra människor.
Fotbollsspelare klädda i gult, blått och vitt uniformer spelar mot andra spelare klädda i guld och blå på en stadion.
Två tjejer tävlar i en motocross race pratandes vid startlinjen.
Tre bicyklister som bär skyddsutrustning medan de tävlar nerför en brant manssluttning.
En person som cyklar i smutsen.
En man med svart hatt, ett par glasögon och ett långt vitt skägg sitter bredvid en målning av sig själv.
En collegestudent tittar på papper i ett rörigt studentrum.
Vid en fullsatt baseballmatch lutar sig slagmannen bakåt och griper tag i slagträet när bollen landar i fångsthandsken.
En kvinnlig artist är barfota och uppträder framför en publik.
En fotbollsspelare ringer en tid ut medan hans lagkamrater förbereder sig för att spela fotboll.
En man som håller i ett stålspö skapar en eld.
En man och en kvinna som bär labbglasögon arbetar med flaskor i ett labb.
Målvakten flyr försvararen för att få bollen till en lagkamrat.
Två lag som spelar mot varandra, ett rött och ett blått med två medlemmar som kväser.
En kemistudent tittar på innehållet när det sitter på en viktskala.
En ung kvinnlig student, som bär en uggla-t-shirt, arbetar med ett experiment genom att fylla sina provrör.
En löpare som bär lila strävar efter mållinjen.
Två män spelar en sport liknande fotboll, med en i rött försöker passera försvararen i blått.
Hjordar av cyklister tävlar av åskådare.
En man i blå uniform hoppar i luften för att skjuta en basketboll.
Promenader och prat och att vända träd till mulch.
Två tonårshonor som flyter på vatten medan de sitter i jättelika plastbollar.
En baseball kanna är att kasta en pitch.
Två män, en med nummer 13 jersey och en med nummer 24, spelar baseball.
En man som spelar gitarr framför en mikrofon.
En man skateboardar i en park, och han är på en vägg, och det finns andra skateboardare i bakgrunden.
En man som står osäkert på en stege och målar en vägg.
En stor grupp människor sitter på en brygga med utsikt över en sjö.
En man som spelade gitarr när han rökte en cigarett.
En grupp människor på isen och en sågade ett hål i den.
Tre barn i havet bredvid en segelbåt.
En äldre man som bär turban sitter på marken medan han håller i en stor sten.
En man i grön skjorta som vinkar medan han går.
Två män, en som dricker en öl, sitter och ler mot kameran.
En tjej i grå t-shirt sitter i en stol.
Det finns en cyklist som cyklar i luften i en utomhusmiljö.
En kvinna på ett apotek tittar igenom en hög med papper.
En man poserar på en skidbräda med snö i bakgrunden.
Vänner visar upp en ny drink.
Ett lyckligt äldre par delar en dans medan en yngre dansande kvinna ser på.
En man poserar bredvid högar av cowboyhattar.
En dansare som bär vit skjorta och shorts fotograferas av en man som också bär vit.
Ett barn tittar genom ett teleskop på en lekplats.
En man tävlar en ovanlig typ av cykel med många människor tittar på honom.
En man som anstränger sig för att avsluta ett lopp
På stranden ligger en man på magen och läser en bok medan en kvinna i en polka-dot bikini solar.
Turister observerar ett geografiskt landmärke genom sökare.
Två cyklister, i gult, tävlar i ett lopp.
Två fotbollsspelare, en i rött och den andra i gult, slåss om en fotbollsboll.
En kvinna med gröna knäskydd åker skridskor inne i ett cementhål.
Det här manliga teamet springer längs grusvägen med kanoten.
Två honor, den ena i mörkblå skjorta och den andra i vit skjorta, spelar lacrosse.
En snöig dag rör ett barn i röd rock vid en dinosauriestaty.
En vit man som utför ett vattenbräde trick i en sjö med träd i bakgrunden.
En kvinna med svart hår och en konstig outfit på.
En pojke med blå kort stå på trafiksignalstången.
Två äldre män bär ytterkläder medan de använder kikare.
En kvinna som bär en grön huvudduk skrattar medan en kvinna i bakgrunden paddlar en båt.
En pojke förbereder sig för att spela basket medan han lyssnar på sin favoritmusik.
En kvinna i svart klänning och hatt rider en enhjuling framför en publik.
En man som håller tal inför en folkmassa.
En umpire och en fångare väntar flitigt på smetens nästa missade boll.
En polis kramar en kvinna på gatan.
En grupp äldre människor som spelar en mängd olika instrument medan de sitter vid ett bord.
Två män som arbetar tillsammans för att rista isskulptur.
En grupp människor, på stranden, en solig dag.
En cricketspelare ställer upp bollen.
En man i jeans overall håller fast vid en hästs leder, som sitter fast i ett dragsystem med en annan häst.
En skäggig man pratar i telefon medan han ser nöjd ut.
Singer Avril Lavigne är hukad på ett knä och håller i en mikrofon.
En skara bicyklister rider längs en gata, med åskådare på båda sidor.
Ett fotbollslag i maroon tröjor tar planen medan hejaklacksledare hejar på dem.
Spelare på fotbollsmatch samlas runt domare som förberedelse för handling.
Två cyklister tävlar i en road race som uppmanas på av publiken som kantar kapplöpningsbanan.
En man leker Frisbee i parken.
Kvinnan håller i en matkasse när flera barn tittar på den.
Två tävlingscyklister rider genom en korridor.
En man på gatan som gör en tavla från ett foto.
Två män som jobbar i en cykelaffär.
Arbetaren koncentrerar sig på sin uppgift som trädgårdsmästare när han pryder häckarna med omsorg.
En kock arbetar hårt när han tar ut mat ur ugnen.
En kvinna spelar för USA volleyboll laget, spika bollen över nätet.
Unga män ser en kvinna gå nerför trapporna.
Fyra män spelar golf på att sätta grönt av ett hål på en solig dag.
Ljusfärgade kajaker som bär två personer vardera paddlas nerför en trädkantad flod.
En man med badmössa och glasögon simmar i en flod.
En man som skjuter en pilbåge mot ett mål.
Färgglada gula platser med en gles publik rad upp bakom fyra fotbollsspelare försöker gå efter en boll.
Snabb cykeltävling i ett främmande land.
En motocross racer i grönt rundar ett hörn och rör upp smuts för publiken.
Cyklare tävlar i en lång blåst uthållighet test.
En cykelförare i ett lopp följs av en polis på en motorcykel.
En kvinna som sjunger in i en mikrofon.
En man i blå hatt och ett förkläde som ristar träfigurer.
En blå restaurang som sitter i vattnet.
En man som sjunger och en man som spelar saxofon på en konsert.
En surfare i luften på sin bräda i havet.
En professionell fotbollsspelare i ljusblått utmanar en annan fotbollsspelare i blå och röda ränder för bollen.
Fem damer klädda i livfulla färger med kul dans.
En cykelförare, i full skyddsutrustning, är upphängd i luften ovanför ett fält av smuts och gräs.
En kvinna med långt hår som går genom en äng
En grupp människor på ett grönt fält hoppar upp och ner.
Smutsig blond man med tatueringar spelar gitarr.
Ett volleybollspel där två pojkar som försöker för bollen, för sitt lag.
En grupp killar satte ihop och roade sig medan de drack.
En cyklist i en vit hjälm rider ovanpå sand vid ett staket.
En baseballspelare, med catcher och umpire visade bakom sig, är på väg att slå bollen.
New York Yankees basebollspelare som slår en baseballplatta.
Folk samlas på en gammal glassbil för att få traditionell glass.
Ett ungt afrikanskt amerikanskt barn som sitter på en gunga med båda armarna som håller fast kedjorna på gungan.
Två tjejer kramas framför en amerikansk flagga.
Bicyklisterna närmade sig vänstersvängen i en flock under loppet.
En blond volleybollspelare når upp till bollen.
Flera fotbollsspelare står på en brun, gräsbevuxen, lantlig åker med en byggnad i bakgrunden.
En man kite surfar i havet.
En flickor volleyboll spel där ett lag bär övervägande vita skjortor och den andra bär gröna skjortor.
En kvinna som slår en volleyboll med två händer.
Två volleybollspelare mot nätet försöker blockera ett skott från det andra laget.
En kvinnlig volleybollspelare ställer in bollen.
En grupp tonårspojkar i gula och blå fotbollsuniformer besprutas med vatten.
En gatuarbetare som bär ljus orange säkerhetsutrustning plockar upp sopor längs gatan.
En vitklädd fotbollsspelare försöker snappa upp en fotboll som snabbt närmar sig målrutan.
En man som sprang på en folkmassarad gata i ett maraton.
En stormästare och studenter i en kampsport klass buga mot varandra i en gest av respekt för varandra och den heliga konsten.
Marathonlöparen Izabella sprang medan de följdes av en skara människor i kostymer.
En scen från ett tävlingsmaraton, inklusive flera deltagare, ner för en crowd-lined city street.
En man kör en vintage racerbil runt banan.
En kvinna i ett hårnät tittar på ett prov under ett mikroskop.
En ung pojke i klänning som blandar färg med udda färgade byxor.
Medlemmar av Baltimore Orioles firar efter en seger.
Fyra fotbollsspelare går över ett fält och håller hjälmarna ovanför huvudet.
En man som sätter på sig shorts i ett rum med några andra människor.
High school fotbollsspelare spooping upp en fumla.
En person som rider på en surfbräda på en stor våg.
En grupp unga män spelar basket utomhus.
Skäggig svart klädd manlig artist visar sin skicklighet genom att svänga en eldlinje i varje hand i bågar.
Gula uniformerade fotbollsspelare som ser sin lagkamrat sparka iväg.
Två fotbollslag, en i gult och vitt, den andra i blått och vitt, spela fotboll.
En man i gul skjorta springer i ett lopp.
Barn, en del i rött och en del i neongult, spelar fotboll.
En hockeyspelare som försöker göra mål
En grupp flickor i blå och vita uniformer är i en cirkel och höjer sina händer.
Veteran rocker utför en hyllning i den dödliga heta solen.
En ung man håller en hammare ovanför en rädd ung man medan en annan vaktar.
Två fotbollsspelare, en klädd i rött och en klädd i blått, spelar fotboll mot varandra.
Det ser ut som om spelaren i bourgogne just sparkade fotboll över # 5 huvud.
En löpare fångas springande mitt i ett lopp.
En liten unge med mat över hela ansiktet i en barnstol.
På den trånga utomhuslokalen, en sångare gester till fansen.
Fyra män spelar fotboll, två i vita tröjor, en i röd tröja och en målvakt i bakgrunden.
Tre kvartsbackar värms upp före matchen.
Två unga stilrena människor går entusiastiskt nerför en stad gata på natten.
En BMX cyklist gör ett stunt på en flodbank över floden från en fabrik.
En svart dam i traditionell klänning med en korg balanserad på huvudet går nerför en strand full av solbadare.
Hockey målvakt i röd tröja redo att blockera ett skott.
Fotbollsspelaren i brun springer med bollen från spelarna i vitt.
Fyra barn i ett låtsasägg som har kul.
En man rider på en motorcykel och blir bevakad av en folkmassa.
En man utför ett trick på en vattenbräda.
En kvinna klädd i en grå skjorta spelar ett hästkapplöpningsspel.
Barn och vuxna rullar skridskor i en skatepark.
En man i jeansjacka och sandaler som fixar sin cykel.
Två män övar dansrörelser medan en dam fotograferar.
Två unga flickor skriver med krita nära en vattensamling.
Det här är en ung kille som sträcker sig efter en falk på en abborre.
En asiatisk man som bär silverpansar över solbrända kläder under sig och håller ett vapen uppe i sin högra hand på en häst som också är prydd med silverpansar.
Jag reparerar taket på en skola vid kusten.
En liten flicka ler när hon bär en vit skål på huvudet.
En man med hattar påsatta i sidled använder en mikrofon.
En man som bär en hustrumisshandlare sjunger in i en mikrofon när ett blått ljus lyser på honom.
Ett antal män rider elefanter genom en lerig flod.
En man i en blå jersey går igenom en baseballmatch.
Folk ser en jockey rida en häst.
En häst och jockey rusar över en flod med en bro full av observatörer i bakgrunden.
En kvinna är på hästryggen, hoppar över en vägg gjord av kvistar och metall.
En rullskridskorska i röda och svarta strumpor och en svart skjorta är armbåga en annan åkare ur vägen.
Band spelar på scenen med Weezer symbol i bakgrunden.
En kvinna formger långsamt en skål med händerna med en lerspinner.
En kameraman filmar en annan man i en grön skjorta på en strand.
En kvinna som bär en brun skjorta tittar genom ett mikroskop medan andra står bredvid henne.
En ung kvinna tittar i ett mikroskop.
En person av asiatisk härkomst bär en blå och svart krigarliknande klädsel, och människor är i bakgrunden.
Två personer tar bilder och tittar på en vacker scen vid vattnet.
Två poliser står på trottoaren när passageraren i bilen tittar på dem.
Man sitter på toppen oljerigg på maskinen fungerar.
Tre personer rider longboards nerför en kulle i fulla läderdräkter och hjälmar.
En grupp människor är på en arbetsbåt som ligger i vattnet.
En grupp på sju personer bär forsränningsutrustning, vit vattenflotte nerför en flod.
Kvinnor på en svängtur på en nöjespark.
En kvinna spelar violin och sjunger samtidigt medan hon sitter i en stol.
En liten flicka borstar tänderna.
Flera män klättrar på en stolpe som en publik tittar på dem.
Två sekreterare samtalar i receptionen på ett hotell.
En ung pojke jagar en fotboll som studsar bort från honom.
En defensiv fotbollsspelare försöker ta itu med en offensiv fotbollsspelare som håller i en fotboll.
En man i grå skjorta lägger glänt till kakel.
En skateboardåkare gör ett trick på en skatepark.
En man vinkar högt i luften, ute i havet.
En löpare sätter hinder över ett hinder.
En ban- och fältidrottare som kör på en röd bana i en stad med många åskådare som tittar.
En idrottsman hoppar över ett hinder.
En manlig cyklist hoppar en ramp i en tävling eller korsar mållinjen.
Tre män arbetar på en cykel, som har placerats upp och ner.
En person, som hukar sig på en surfbräda, surfar i en vattenförekomst.
En man i blå uniform som jobbar med mekanik.
En mörkhårig pojke med en grön t-shirt spelar i en vattenfontän medan två andra tittar på honom.
Flera arbetare står på och runt en stege.
Tre män med hårda hattar och säkerhetsanordningar sitter på en båt och en bro är i bakgrunden.
Barn i klassrum med uppstoppade djur.
2 personer engagerade i samuraj stil strid i en gymnastiksal.
En man som njuter av dagen vid vattnet och väntar på att få dela ut ballonger.
En kvinna i svart skjorta sitter framför ett mycket stort konstverk i ett stort rum.
En mountainbikeer hoppar över ett hinder.
En man står upp och snurrar ett lerkärl på sitt lerkärlshjul.
En svart man står utanför ett museum och pekar på det.
En domare höjer handen på en brottare som bär grönt medan en brottare som bär blått ser på.
Två tjejer i bikini som spelar volleyboll på stranden
En liten grön bil med nummer 63 på dörrkapplöpningarna på en kärrväg.
Två män i skyddsutrustning sågar genom metall.
Militärer i vita uniformer står sida vid sida.
En tjänsteman konsulterar en konkurrent vid ett kampsportevenemang.
På den här bilden kör två tjejer karate.
En liten pojke i jeans, röd randig skjorta och sneakers, sittande på trädgrenen.
En kvinna i svart skjorta och khakibyxor sitter på golvet och drar på bruna högklackade stövlar över rosa och röda strumpor med hjärtan på.
En gammal man syr kläder på en trottoar.
En man klädd i en långärmad, knäppt blå skjorta och en svart och silverfärgad keps håller en telefon i örat.
En racer firar sin seger genom att hålla är trofé och duschas av champagne.
En hund hoppar högt upp i luften i landet.
Orange motorcykel racing runt en böj i ett racetrack.
En person placerar okokta hamburgare pattys på en kolgrill.
En man med glasögon som håller i en statys svans.
En publik hejar och passerar streamers på en stadion medan en blå flagga vågor.
Två kvinnor klädda i svart lutar sig bakåt på vita bord.
Under en rugbymatch tävlar spelare från båda sidor om den lösa bollen som lagkamrater tittar på.
En kille med svart hjälm, rider mountainbike.
En man försöker åka skidor på den sista snöplätten som finns kvar på kullen.
Två personer bär hjälm och solglasögon en solig dag.
En liten pojke klättrar på apbarerna på en lekplats.
En man står i en kyrka medan folk runt omkring honom tittar.
En man klättrar uppför en klippa med en skog i bakgrunden.
En mor hjälper sin dotter att klä sig för ett speciellt tillfälle
Tre personer på cyklar på en smutsig kulle, en är i luften.
Två pojkar hoppar och får luft över en ravin med mountainbikes.
Två män sitter på en vit soffa i ett vitt rum med separata bärbara datorer.
Två bilar som är inblandade i racing kör mycket nära.
Fotbollsspelare på ett fält med en boll som går in i nätet.
En man som åker skateboard uppför en lutande ramp.
En man i beigedräkt sitter vid ett träbord med fem barn och ritar bilder.
Två personer tävlar i en fäktningstävling.
En äldre man med skägg i mörk kostym går genom en regnig stad.
En kvinna med kort blont hår försöker fixa sitt hår
En bebis tuggar på fingrarna medan han bär en blå randig klädsel.
Den lokala elektriska arbetaren hänger upp några ledningar.
En ung blondhårig man skrattar när han tar av sig skjortan i en offentlig miljö när åskådare tittar på.
En kvinna använder en ostgröt.
Två män står på en medelstor fiskebåt i havet, när solen går ner bakom dem.
Fem barn är på en fotbollsplan på väg mot målet.
En man i gul overall står på ett podi och tar emot en trofé bredvid en man i rött och med overall.
Ett ljust klädd barn går i en sjö.
Ung punkrock gitarrist, bär en röd fodrad jacka med en bricka, är framför dimmig blå och lila belysning.
En man som gör ballong och njuter.
En ung man sprängde ballonger för att tillverka djur åt de sju upphetsade barnen som såg på.
En äldre kvinna använder ett spinnhjul för att skapa tyg.
En man tar på sig rollen som återförsäljare och sitter vid ett kortbord.
En liten flicka i lila hatt som sitter under en kundvagn i en livsmedelsbutik.
Fem små barn är engagerade i en fotbollsmatch.
Två personer är på en båt i vatten.
En man som cyklar på ett fält.
En man går över en fotbollsplan klädd i rött och vitt.
Televisionskameror för att spela in en jämn på en teater.
Ett barn får sina tänder borstade.
Två män klädda i Red Bull varor firar genom att öppna drinkar tillsammans vid ett evenemang.
En man och en kvinna som håller hand framför en sjö.
En person som bär våtdräkt rider en jetski in i en våg.
Tre killar i röda uniformer firar ett mål i en fotbollsmatch.
En man i en röd hjälm rullskridskor nära stranden med två hundar i koppel.
En man som driver en jetski gör en volt i vattnet, och ses upp och ner.
En person, i ett kök, håller ett ägg ovanpå en skål med ris i.
Fyra unga pojkar som spelar fotboll och jagar en vit och röd fotboll.
En man och en kvinna som ler medan de ser på när någon gör creme brulee efterrätt framför dem.
En person i SCUBA-utrustning står framför ett vidsträckt vattenbredband.
En blond tjej som bär en svart och vit boa poserar för kameran på en mycket trång plats.
En pojke lutar sig mot en tegelvägg nära några träd.
En man som rider en röd och vit cykel på solig dag.
En äldre man sköter om en trädgård.
En forskare i en labbrock använder ett mikroskop.
En grupp flickor står på en fotbollsplan och poserar för kameran.
En man klädd i svart och guld över rock rider en svart och vit häst.
En del fotbollsspelare vid sidan om tittar på när en lagkamrat börjar spela.
En fotbollsspelare förbereder sig för att kasta fotbollen när resten av hans lag klockor.
RollerSkaters slåss ut på betongen.
Två lag män, ett lag i blått och det andra i kamouflageuniform åker skridskor.
Två personer tävlar i ett motorcykellopp.
En äldre herre som försöker reparera en uppochnedvänd cykel nästa också ett silver fordon.
En flickas volleyboll lag har en match.
Den vackra damen i vitt dansar balett framför en stor, vacker fontän.
Ungt kvinnligt volleybolllag står vid sidan om för att förbereda sig.
Vacker dansare i röd kjol och hon slår en pose med benen i luften.
Tre barn skriver uppmärksamt i ett klassrum.
Två kvinnor sitter på en svart soffa med kläder och en handväska däremellan.
Ett par som står ute och omfamnar och tittar över landet.
Några personer står i ett klassrum längst bak i rummet medan man sitter vid ett skrivbord.
Två kvinnor beundrar hängbron från sidan.
En fotbollsspelare försöker tackla en spelare i motståndarlaget som kör med bollen.
2 unga pojkar i pisswee fotbollsmatch
En ung rödhårig kvinna letar efter mål på skjutbanan.
En Ohio State team maskot utför på fältet.
Två små barn en pojke och flicka färglägger vid bordet med sina crayola kritor och lite papper.
En segelbåt med många människor seglar på vatten.
En man i en grön jersey och rullskridskor snubblar när en man i en svart jersey verkar kollidera med honom.
Två små barn klädda som Spider Man åker nerför en rutschbana.
En kvinnlig simmare kommer upp för luft som hon gör fjärilen stroke.
En grupp kvinnliga simmare dyker ner i en simbassäng.
Fotojournalist på en motorcykel, följer maratonlöpare, en bär en grön skjorta och skor, den andra fluorescerande orange med blå skor.
En mycket vältränad kvinna löper med bladverk i bakgrunden.
En artist hoppar från scenen in i en massa fans.
Två personer, en man och en kvinna, sitter utanför.
En dam i röd skjorta med rött hår skrattar medan hon kastar en kudde över sin vänstra axel.
En ung man i grön och vit randig skjorta som spelar rullskridskohockey.
En man i orange och vitt rider sin mountainbike genom en skog.
En röd ekorre på en trädgren med gula blad i bakgrunden.
Ett barn tittar genom ett mikroskop medan vuxen står vid kanten av ett bord.
Ett par, klädda i svart, vinröda och vita, dans.
Ett militärt kirurgteam, ett i kamouflage, utför en operation på ett fältsjukhus.
Två lag, ett med svarta uniformer och ett med blå randiga uniformer springer nerför en idrottsplan.
En liten pojke med brunt hår och en tröja ler busigt av några blommor och växter.
En kvinna som bär en blå kjol är på en gångväg och tittar på en vattenförekomst.
En fotbollsceremoni i en fullsatt stadion med laget som förbereder sig för att buga och ta bilder.
Två idrottare fäktas i en fäktningstävling.
Två män slåss mot varandra i fäktning.
Två personer stängsel och en förlorar sin sko.
En man i bruna byxor och en randig t-shirt som jonglerar med tre vita nålar.
En manlig labbarbetare med glasögon undersöker något med hjälp av ett mikroskop.
En vattenpolo händelse äger rum med en gul boll i en pool.
En pojke som bär skyddsglasögon använder ett lödjärn på en elektronikbit.
En person på en cykel rider på en grusväg i skogen.
En manlig snowboardåkare fångar lite luft och gör ett trick.
Ett barn leker på stranden och stänker vatten överallt.
En kvinna är på ett gym och tränar på ett löpband.
En man lyfter upp en kvinna i rosa klänning under en dans på en föreställning.
En fotograf som fångar en skateboardåkare mitt i tricket.
En ung pojke med blått hår och stora blå ögon borstar tänderna
En grupp människor står på en rörlig trottoar.
Redo och ställa som två hockeyspelare på isen vänta med pinnar ut framför dem, förutse pucken.
Människorna verkar uppskatta pojkarnas ansträngningar på scenen.
En kastare har precis kastat bollen mot smeten på ett baseballfält.
En basebollkastare kastar en boll.
Två män poserar för en bild medan de förbereder sig för att ta en drink.
En baseballspelare kastar en tonhöjd från högen.
En svart, röd och vit tävlingsbil zoomar förbi på en grå bana med en blå kant, skarpt i fokus jämfört med en suddig publik i förgrunden.
Folk äter på en restaurang, en del äter medan andra beställer.
En kvinna och en ung man som skrattar i ett sovrum.
En näsduksklädd man sopar skräp vid en händelse.
En fotbollsmatch för pojkar äger rum, och en pojke i en vit tröja sparkar bollen.
En man blåser in i en lång pipa
Det finns två kilted män, en av dem äldre och håller säckpipa med den andra med en trumma.
En grupp män som bär kilts kastar en lång träpinne.
En man i svart skjorta och grön rutig kilt kastar ett långt träspjut, som flera män tittar på från sidlinjen.
En kvinna i orientaliska kläder poserar på en grön matta.
Flera män cyklar nerför en hall i ett evenemang på en solig dag.
Folk som cyklar i ett lopp.
En racerbil går förbi på racerbanan.
En cyklist driver hårt för att slutföra ett lopp.
Två simmare i vattnet, var och en i sin egen fil, samlar ett andetag mitt i slagfältet.
En man som sopar trapporna ner från sitt hus.
En ung vit man med svart hår, svarta byxor, och en vit och svart polka-nedsatt skjorta håller och sjunger in i en mikrofon.
En gymnast bär en livvakt och gör ett handstånd.
En tennisspelare slår en tennisboll med all sin kraft.
Marathonlöparen fokuserade på löpningen.
En grupp kvinnor tävlar.
En vit, manlig, professionell cyklist rider på landsbygden.
En kvinna som sitter på en tygbit omgiven av smuts och arbetar på en tygbit
Tre manliga vänner i shorts står tillsammans och pratar.
En föreställning sätts på av många flickor i vitt.
En maratonlöpare joggar förbi fotgängare och bärbara toaletter.
En ung vuxen läser en bok på tvättomaten medan han väntar på att hans tvätt skall göras.
Kenyanska kvinnor springer i ett maraton.
En man som bär hatt är skateboard framför en graffititäckt vägg.
Flera kvinnor springer i ett lopp, medan publiken tittar på.
Houston Texans quarterback håller en fotboll mot Minnesota Vikings medan hans running back rör sig mot bollen.
Två fotbollsdomare väntar på bänkar med träd i bakgrunden.
En fotbollstränare med vit skjorta och svart visir har armen runt en av sina spelare på sidlinjen.
Två spelare möter varandra under en fotbollsmatch nattetid.
En man i blå baddräkt hoppar från en klippa ner i vattnet medan en annan man tittar.
Barnet sitter på klipporna vid parken.
Två män boxas i en boxningsmatch i en ring den ena har röda shorts den andra har vita shorts båda i kampen stanza.
Det röda laget jagar bollen under flickornas fotbollsmatch.
Kvinna i blå shorts och vit skjorta sparkar en fotboll.
Ett par kysser varandra medan någon fotograferar dem.
En kvinna i grön skjorta som håller en cigarett särar armarna i en gest.
De tre landhockeyspelare klädda i orange gör för bollen.
En man i hätta knäböjer och böjer sig framåt för att undersöka en motorsåg.
Grupp av ballerinor i vit tutus gör dig redo att dansa
Aggressiva åtgärder händer av målet i denna hockeymatch.
Två personer spelar vattenvolleyboll och en lagkamrat slåss mot en annan.
I köket i en tjusig restaurang har en fin maträtt tillagats av personalen.
En kvinna som säljer mat vid vägkanten.
Två kvinnor tävlar i kampsport evenemang på ett gym.
Två killar i karateuniform sparrar på en vadderad matta.
En kvinna bär en röd se genom tyg över huvudet.
Flera människor går längs trottoaren och transporterar saker till sin nästa destination.
En flicka som bär blå byxor och en skjorta med huva ses flyga upp över nästan två meter från marken och hålla ett glas som hon har tagit bort från diskmaskinen.
En kvinna med hink som städar en offentlig sittgrupp.
En pojke kastar ett föremål framför en glasbyggnad.
En man i en kajak vilar ovanpå en dykbräda.
En ung man i sina boxare gör ett roligt ansikte och sätter på sig jeansen.
En äldre man hoppar fallskärm.
Två män spelar hockey, med en på marken och den andra sprutar honom med is.
Mr Soccer-spelare i det gröna laget försöker skjuta.
En man i blått, som håller två fiskestolpar med den ena pekande uppåt och den andra i vattnet med fisk fångas.
En kvinna hoppar i luften på en trädfodrad stig på en höstdag.
Tre män spelar fotboll där en kille bär röd uniform håller i fotbollen, den andra killen bär röd uniform och den tredje killen bär vit uniform.
En Texas A&amp;M fotbollsspelare som kör med bollen.
Det finns en grupp av nio unga kvinnor som bär långa svarta klänningar med mappar, står på metall blekare och sjunger inför en grupp människor.
De här två männen ska ta bollen på en fotbollsmatch.
En man i klänning dansar när en annan man står vid en stege och vänder sig åt andra hållet.
Texas A&amp;M: s Ryan Tannehill är nästan sparkad av en Iowa State spelare.
En korsvakt hjälper folk att ta sig över gatan.
En husky kvinna med röd hatt, styr trafiken.
En man i blått med munnen öppen bredvid en medicinsk apparat.
En gammal man som svettas håller ansiktet i handen.
Några män springer maraton med folk som hejar på dem.
En kvinna på en cykel racing.
En medelålders man är förfärad eftersom någon vill att han ska prova en spett med några udda fiskar på den.
En man tränar utomhus.
Ett fotbollslags spelare i den blå och guld uniform kör ner 30 yard linjen mot slutzonen.
En man klädd i rosa rider en cykel i ett lopp.
En kvinna som bär vitt drar av ostblock från en transportör.
Mannen i röd skjorta lyfts av sina lagkamrater.
En vit pojke i gul och afrikansk-amerikansk flicka i lila är av orange skåp.
Flera män i gröna och röda uniformer spelar fotboll.
En kvinna cyklar i förgrunden med andra cyklister i bakgrunden.
Människan är fast besluten att cykla sin väg till mål!
University of Iowas Hawkeyes fotbollslag, gör mål i slutzonen mot Michigan State Spartans.
En mycket söt ringbärare kysss motvilligt av blomsterflickan.
En svart flicka i lila jacka tittar på en bok, när hon sitter på en färgglad stol.
Två fotbollsspelare faller till marken nära bollen.
En svart och vit hund hoppar upp ur vattnet och en brun hund skakar av sig.
En man, som går sin pommern, ger en cyklist vägbeskrivning.
En middagsbjudning äger rum med många människor som alla bär kronor och äter mat i en ljust upplyst matsal.
En proffscyklist i blå, gula och vita cykelkläder.
Två honor befinner sig i ett kemiklassrum; en häller en lösning i en bägare.
Förhoppningsvis har jag ögonbryn när jag blandar dem.
En grupp unga gymnasieelever ler medan de utför ett vetenskapligt experiment med bägare och överföring av vätskor
En vetenskapsman som är djupt inne i sitt experiment.
En stor kvinna med rosa fjäderboa promenerar nerför trottoaren.
En man klättrar en stenblock över en vattensamling.
Tröjalös ung man som klättrar uppför klippan och letar efter nästa handtag.
En man bär många stora väskor som är fastsatta på en stolpe.
En manlig löpare i en orange och vit t-shirt och svarta shorts sprintar längs banan.
En ung man som fick medalj och hängdes runt halsen.
En person i en regnbågsfärgad snödräkt åker snowboard nerför en snöig sluttning.
En man som sjunger och spelar akustisk gitarr i ett offentligt område.
Tre cricketspelare är i aktion på ett mycket grönt fält med palmer i bakgrunden.
Två män i svart firar på en tennisbana mittemot två män i vitt.
En ung kvinna sitter framför sin dator och försöker studera det finstilta på ett papper med hjälp av en läkares spotlight fäst vid hennes huvud.
Lärare framför klassen som läser en bok högt för grundskolebarn.
Tre personer står med fiskestolpar på klipporna nära vattnet.
En man som bär jersey nummer 39 spelar hockey.
En grupp människor tar bilder på en gångväg framför en stor vattenförekomst.
En löpare stänker genom en stor pöl i skogen.
Två män sitter på toppen av en väderskadad fortliknande struktur bredvid havet, fiske.
En pojke spelar fotboll på en lekplats.
En kille utan tröja klättrar upp för en sten.
Två män försöker ställa in sitt teleskop som är placerat i ett fält.
En ung asiatisk pojke, som bär pyjamas, sitter på golvet vid sängen och tittar på en insekt gjord av legos.
En händelse äger rum i ett japanskt tempel.
En basketspelare hänger i en basketkorg vid fötterna, skrattar och pratar med en domare framför en publik.
En man som är vattenskidare och plaskas av vattnet.
Den här mannen i kajaken tycker att kajaken är alldeles för liten för honom.
Arbetare flyttar tegelstenar från en vit och grön lastbil.
En liten tegel gränd med en man som går i slutet
En skjortlös man ligger på gatan.
En kvinnlig simmare med goggles och en mössa gör backstroke.
Aaron Rodgers ler mot Donald Driver som står i slutzonen.
En man klädd i sportutrustning och solglasögon sitter i en båt, paddling med en stor åra.
En ung man på gatan som gör ett skateboardtrick.
En leende flicka bär en Speedo baddräkt, glasögon och mössa med händerna på pannan.
Fyra damer och en man som övar musik i ett vardagsrum.
En blond kvinna går framför en grupp på tre personer.
En blond tennisspelare i aktion på en gräsbana.
Två personer arbetar på ett kafé
En kvinna läser en tidning på tunnelbanan.
En person fångar en våg på en surfbräda i havet en klar solig dag.
Två pojkar leker med stora pinnar på gården.
En man som går på brädor medan han håller fast vid en stor stege lutar sig mot ett hus.
En man försöker ta tag i sin stege stående på byggnadsställningar.
Latino man håller skylt på trottoaren utanför främja Quiznos-Subs.
Ett manligt och kvinnligt team av rullskridskor är i kostym och uppträder i en tävling.
En man läser tidningen på ett däck under några träd.
En cyklist på neongul cykel är luftburen.
En dirt-bike racer tar en hård sväng på en smutsbana med en åskådare i bakgrunden.
En man kör en liten motorcykel genom en upptagen marknad.
En man som bär gula leenden mot kameran när han står med en kalkon som kommer ut ur ugnen.
Panelrepresentanter som sitter på en scen i en auditorium.
En grupp människor i gula och svarta uniformer uppträder framför en stor publik.
En demonstration mitt på en fullsatt flygplats.
En liten flicka i en vit solklänning ler och glider ner för en blå rutschkana.
En man och en hund leker dragkamp.
Fyra unga pojkar ställer upp sig vid startlinjen för att köra ett lopp
En grupp kvinnliga idrottare är sammanflätade och upphetsade.
En kvinna matar en äldre man med tårta vid en bröllopsfest.
En sen kvällsmatstånd tar kundernas order.
Tjejen i köket blandar smet i en skål för våfflor.
En man som skateboardar på gatan med upplyfta armar.
En hane i vit t-shirt och denim shorts skateboard nerför en stig.
En kvinna med röd skjorta och glasögon driver en orange övning.
En mountainbike racer på en grusväg under ett lopp
Den här mannen jobbar med en I-pad.
En brun hund och en vit hund springer över en stenig kulle.
Tre unga män spelar fotboll på stranden i shorts och strandkläder medan vissa människor tittar
Ett blått lag och ett vitt lag tävlar om att vinna ett sportspel.
En man i svart skjorta och en brunhårig kvinna som sniffar flaskans innehåll.
En grupp människor står och äter som en man i en vit jacka och pekar finger.
En grupp människor som spelar musik offentligt på unika instrument.
En basketspelare förbereder sig för att kasta bollen i ett spel på skolans gym.
En person som bär en rosa skjorta och cyklar på en grusstig.
Tre mariachibandsmedlemmar spelar på en gräsgård.
En byggnadsarbetare hjälper till att anpassa cementplattan på vägen.
En liten brunhårig flicka uppe i ett träd.
En person på en cykel hoppar över en gruskulle.
En ung pojke på rullskridskor hoppar över en blå tunna.
Barnen med julhattar dansar glatt runt julgranen.
En snowboardåkare slipar på en räls i ett snöigt, bergigt område.
Tre personer, två män och en kvinna rider i en båt.
En förare i racingutrustning och en hjälm kör en elegant, blå motorcykel.
En man på en gul och grön surfbräda nära stranden.
En man som hamrar en spik på en träbit i bara fötter.
Två forskare undersöker ett mikroskop omgivet av komplexa maskiner.
En man med långt lockigt hår som grymtar som en man använder en klippare i skägget.
Män borstar is för att flytta vikten till målet.
En grupp dykare räddar en man i vattnet.
Två personer njuter av en praxis av en oidentifierad glidspel.
Tre personer på en hockeyring spelar någon form av spel.
En man med en gulgrön tröja som sparkar en fotboll.
En grupp unga män klädda i lila förbereder sig för att fånga en lagkamrat.
En kanna står vid högen och kastar.
En man, i mitten av swingen, spelar cricket med en komplett cricket uniform på en idrottsklubb.
En liten flicka får hjälp med sina leksaker.
En person i en tomtedräkt hälsar på barn utanför en byggnad medan föräldrarna tittar på.
Två seniorer och en kvinna dukade ett bord.
En ljusblå tröja idrottsman gör sig redo att ta emot passet mitt i hans grå skjorta motståndare.
En kvinna springer ett maraton i en park.
En man rider en BMX cykel med en skog i bakgrunden.
En cyklist cyklar i skogen.
Medan man spelar fotboll, börjar en man i gult falla, medan en man i vitt snubblar över honom och trampar på sin fotled i processen.
Man poserar för en bild med sin flickvän.
En basketspelare klädd i vitt tittar på sin motståndare, som är klädd i svart, dribbla en basketboll ner på banan under ett spel med åskådare.
En person rullskridskor med knäskydd, hjälm och handledsskydd.
En tjej med nummer 3 på tröjan går över ett gymnastikgolv.
Två ungdomar deltar i en vänlig snöbollsmatch.
En man ligger bredvid en flod och röker en cigarett.
Mannen klädd i löparkläder går längs gatan.
Båt på vattnet i Wien rodes av män med randiga skjortor.
En man sover utomhus med sin bokväska som kudde.
En man med vit skjorta och blå shorts lutar sig över en kanot i slutet av en docka.
En grupp människor som står över ett bord.
Ett yngre par som sitter nära varandra samtidigt som de njuter av en 3D-film.
Kommentatorer och programföretag där både i en arena före matchen.
Penn State basketspelare, nummer 11 skjuta för korgen med bollen bara lämnar fingertopparna.
En person med kort blont hår och glasögon ser förvirrad ut, medan han står framför många porträtt.
Två lag av män spelar basket på en bana i en tom stadion.
5 basketspelare försöker få bollen.
Basketspelare som spelar inför en liten publik
En kvinna och ett barn sitter på en stock och tvättar kläder.
En ung pojke sitter på en strand och fyller en vattenflaska med sand.
Två barn leker Jenga på ett trägolv.
En man utför kampsporter på en annan man i ett gymnasium.
En kvartsback passerar en fotboll under en NFL-match.
Skateboarder hoppar från en fem meter hög klippa och utför ett stunt.
En mc fixar däcket på en solig dag.
Två kvinnor med svarta klänningar och röda toppar står bredvid ett staket leende.
Två damer, sedd bakifrån, en tittar genom ett myntstyrt teleskop
Åskådare sitter i publiken på en hockeymatch medan en fotograf tar bilder från en låda mellan de motsatta lagen.
Föreställare i ljusa kostymer och masker står inför en asiatisk publik.
En person i svarta och vita kläder och en mask är i förgrunden för en grupp barn.
En ensam man sitter i en hamn och spelar dragspel.
En ung flicka, som bär sin laguniform, förbereder sig för att slå en boll, när en annan flicka tittar på.
En man som aktivt surfar på en våg.
En surfare i våtdräkt fångar en fin våg att rida på.
En man som snowboardar nerför en kulle.
En man som rider en blå jetskida är luftburen efter att ha gått över en våg i havet.
Två svarta och vita hundar leker tillsammans utanför.
Två mycket små barn, med färgmärken på sig, målar en mycket röd och gul duk.
En man som rider på en svart snowboard hoppar när folk i bakgrunden tittar på.
En man i grön skjorta och svarta shorts har hoppat upp i luften och är på väg att kasta en röd och vit boll.
Två unga män i en kampsport ring deltar för en publik.
En asiatisk kickboxare är mitt uppe i att sparka sin motståndare i ringen på ett Mohegan Sun casino.
Fem fotografer fotograferar medan en arbetar på sin utrustning.
En ung snowboardåkare fångar lite luft på sin svarta snowboard.
En grupp män som spelar utomhussport.
En gymnast balanserar mellan två räcken med en arm och hans ben är i luften.
Två män, en klädd i blå skjorta och byxor och en klädd i lila skjorta och svarta byxor skapar keramik.
En ung kvinna som spelar gitarr och sjunger på en scen.
En surfare i våtdräkt rider en våg.
En kvinna klädd i svart och en man klädd i vitt trycker på en soptunna.
En man som står i bergen och håller i en pistol.
En asiatisk man i jacka, glasögon och sandaler är på hög höjd och siktar på en pistol.
En tjej med brunt hår som sätter upp ett ljus för en show.
En ung flicka i baddräkt och glasögon sitter och väntar.
Tre män samtalar på en bänk i ett museum.
En man och en kvinna står bredvid skulpturer och pratar medan en annan man tittar på andra skulpturer.
En fotbollsspelare som bär svart försöker ta sig an en fotbollsspelare som bär vitt.
En gammal gentleman spelar musik på gatan för pengar med en ung pojke vid sin sida.
Fyra arbetare i hårda hattar står tillsammans på en arbetsplats.
Tre flickor hoppar upp i luften med uttryck av spänning.
Två kvinnor står i ett kök och torkar ner brickor
Det finns fyra barn som övar vad som verkar vara karate.
En kille som håller tvätten mot väggen medan han pratar på mobilen.
Två fotbollslag på ett fält ett lag klädd i blått en vit den andra klädd i vitt och blått.
Två killar äter en lunch med smörgåsar och chips.
Man med grön hatt och vit skjorta med te med en man i svart huva jacka och glasögon.
En man i hatt och ett förkläde jobbar på en cykel.
En ung flicka i baddräkt gör sig redo att tävla.
En ryttare står för ett ögonblick ovanför sin dirkcykel.
En man ligger i snön medan en flicka står bredvid honom.
En ung man dunkar en basketboll.
En afrikansk amerikan som snider bilder till en planka av trä.
5 barn japaner med bågar tränar framför sensei.
En grupp kaukasiska människor sjunger och håller i musikböcker för att vägleda dem.
Indiska kvinnor spelar musikstolar med vit kvinna.
Två manliga musiker på scenen, klädda i t-shirts och en spelar gitarr, den andra sjunger.
En orkester spelar på en utomhusplats.
Ett gäng barn i ett klassrum som inte gör något arbete.
Folk samlas för ett bröllop.
En kvinna som kysser kinden på en ung pojke i en svart ärmlös t-shirt.
En ung dam som ler i en pool.
Intensiteten i ett ögonblick under en ishockeymatch.
Två män spelar professionell hockey
En kvinna som bär bikini simmar under vattnet.
En ung pojke som äter chokladglass med en sked.
Barn i ett klassrum står uppställda med händerna på varandras ryggar och bildar ett tåg.
En leende kvinna i rött poper korken på en flaska med en pojke tittar på.
En liten flicka är på en lekplats gunga medan en rödhårig man i en grön tröja står förbi.
En kvinna med vit blus får ett porträtt gjort av henne.
En flicka pekar på en plats på en karta i en park.
En tjej i baddräkt, badmössa och glasögon.
En familj tittar ut genom ett fönster och tittar på folk som håller parasoller i dagsljus.
Två män framför musik på gatan framför en tegelbyggnad.
En man med flätat hår och skägg står framför en byggnad och pratar eller sjunger in i en mikrofon.
En kyrkokör framför en julsång medan en projektor i bakgrunden visar texterna.
En volleybollmatch och en man i gul och blå uniform spetsade bollen över nätet förbi tre försvarare i röda uniformer.
Två unga män springer genom gräset på hösten.
En liten flicka kramar en kattunge medan hon tittar på julklappar och en äldre kvinna tittar på.
En person som bär en blå skjorta och khaki byxor klättrar i ett träd.
Tittar genom fönstret i en asiatisk frisör butik medan några kunder har sin frisyr.
En handbollsspelare förbereder sig för att kasta i ett hav av försvarare.
En man i en röd tröja skateboard medan en man i en blå tröja filmar honom.
Köparna letar efter julklappar på Harrods varuhus.
En kvinna i svart baddräkt håller fast vid kanten av en pool.
En kvinna i baddräkt går ut genom en pool.
Fyra kvinnor sitter på gröna utemöbler på en uteplats med ett litet hundhus i bakgrunden.
En skara ungdomar sitter på gräset.
Vuxna och barn njuter av poolen, en del är i poolen och en del sitter runt poolen i solstolar.
Grupp av män börjar en fot ras.
En äldre man spelar gitarr på en rullstol på en stadsgata.
Två poliser sitter på en ohyggligt gul motorcykel.
En man och en kvinna klädd i halvformell klädsel visar ansikten av spänning tittar över ett bord med Jenga block utspridda över det.
En fotbollsgrupp i grön och vit klänning med en gruppbild tagen.
Som målvakt i en gul jersey ser upp i fjärran, en spelare från motståndarlaget i en grön jersey på händerna och knäna har hans ansikte i gräset.
Två musiker spelar musik i en lada.
Ett barn på en torg stirrar ut några stora flytande bubblor.
Kvinnlig besökare som läser karta som beskriver den vattenväg som står framför henne.
En svarthårig kvinna använder sin sminkborste på en annan kvinna medan hon håller upp lillfingret.
En brud håller sin bukett och tittar tillbaka på folkmassan.
En brud med en bukett blommor står bredvid en man i en smoking.
En brud kliver ur sin bil i sin vita bröllopsklänning.
En BMX cykelförare i röda kläder och en hjälm rider sin cykel bredvid ett trästaket.
Ett band spelar medan publiken tittar på dem på scenen.
En ung flicka i blå byxor och en flerfärgad randig skjorta hoppar i luften.
En lärare och hennes assistent hjälper en grupp småbarn med sång eller träning.
Det finns två barn klädda i sina vita karatedräkter, som står och tittar på något eller någon.
Fyra personer står i vattnet och tittar på en jetski, medan en man fiskar i närheten.
En person på en cykel täckt av lera från topp till tå.
En skidåkare går nerför en sluttning.
Ett leende barn sitter i en vit baby utkastare omgiven av leksaker.
En trio av musiker som spelar på en bar.
Pojken i grått tar bilder på sin vän i den randiga tröjan och gör tricks på skateboarden.
En ung man utför ett skateboard trick över några trappor.
En man i blå skjorta som fixar en cykel i ett gult rum.
En hund hoppar för att fånga en röd boll utanför.
En svart och brun hund med en röd boll ovanför spelar i gräset.
En liten hund försöker fånga en röd boll.
Två leriga idrottare från motsatta lag går huvudet till huvudet i en omgång rugby medan fans tittar förväntansfullt.
Två personer Kayaking på det stora öppna vattnet.
Ett barn som bär halmhatt med ett blått band som dricker ur en rosa kopp.
På hörnet hittar du en dam som sitter på sina väskor och sprutar kronan med vatten när de går förbi.
En ung kvinna hoppar så högt hon kan för att bevisa en poäng för sina vänner.
Ett barn i röd rock i ett snö fort.
En liten hund springer bakom en röd boll kastad mot buskar.
Mannen ger den andra mannen en frisyr.
En man i svart tröja och röd skjorta spelar trumpet vid ett träd.
En ung man utför ett hopp på en skateboard medan en annan ung man fotograferar sitt stunt.
En man står mitt i scenen med en mikrofon när lågor skjuter uppåt bakom honom.
Två hockeyspelare slåss över ett mål med hjälp av sina puckar på isen mark.
En man i hård hatt arbetar nära en container.
En man i en mörkblå bil kör förbi några förvaringsvagnar.
En medelålders manlig snickare använder en borrpress i en fullsatt verkstad.
En äldre man i en verkstad bär glasögon.
En glad asiatisk familj poserar för en semesterbild framför den öppna spisen.
Det finns tre barn i sportuniform på en fotbollsplan.
Konkurrerande flickor volleybollspelare försöker kontrollera bollen i luften.
En man står på ett fält med en grön växt i sig.
En man står utanför för sig själv bredvid några gamla byggnader och en tegelgata.
Män klädda i rött och vitt spelar musikinstrument.
En grupp människor som bär blå och vita diskadorhar alla ridande orange cyklar.
En person som leker med en sten bredvid lite smutsigt vatten.
Någon klädd som tomten, fru Claus, och två andra människor rider i tomtens släde, dragen av en häst, genom en snötäckt stad.
Killen i jeans skateboard mitt i natten ett lager.
Två personer går parasailing på havet med en vacker naturskön utsikt i bakgrunden.
Person som parasailing med en styrelse i havet.
Tre män som bär vita skjortor åker skateboard på en väg medan en man och en kvinna tar bilder från båda sidor av vägen.
En DJ med solglasögon och en röd skjorta spelar musik.
En äldre man sitter och tittar på sin datorskärm med ansiktet i händerna.
Man på snöskoter avfyrar upp i luften.
Flera personer i svettkläder låg tillsammans på ett gymnastikgolv, medan en stående person tar tag i ett av sina ben.
En kvinna som bär en blå och gul kroppsdräkt rider en gul cykel.
En cyklist på sin cykel bär en orange och blå kostym reklam Rabobank.
Små barn tittar på en tågsätt som är placerad inom grönska.
Gula, röda och blå flaggor flyger i himlen när en dykare sträcker sig helt i luften.
En manlig gatuartist som går en lina.
En man i svarta oxfords, jeans och en lagergrön över svart skjorta hoppar framför en nedsliten industribyggnad.
En man och kvinna i ett kök med plastmuggar med vin eller champagne.
Två personer i vinterkläder och en hund går längs en strand
En kille som surfar i havet.
Simma ner i vatten utför en flip medan flera kvinnor i bakgrunden titta på.
Tre män har platser första, andra och tredje i ett evenemang och står på podier.
Tre unga flickor tittar på en skärm som en av dem pekar på skärmen.
En man som spelar pingis medan ett barn tittar.
En man med orange shorts och en blå mössa är i ett träd.
Tre hockeyspelare i röda tröjor står tillsammans och håller hockeypinnar.
En kvinna i svarta byxor och en vit skjorta är bergsklättring.
En grupp unga män samlas under ett träd.
En äldre kvinna med glasögon serverar sig själv Raclette i ett rustikt rum.
Tre barn övar karate.
Två personer i gul kajak kommer mot en större vit kajak på öppet vatten.
En asiatisk kvinna klipper en annan kvinnas hår
En kaukasisk kvinnlig frisör klipper håret på en ung vit man som bär ett svart gardinomslag.
En ung kvinna ritar bilder på en vit yta.
En man med mikrofon och två tonåringar studerar något i sina händer.
En man som klipper hår.
En kvinna i en grön topp lyfter en metallskål från spisen.
En grupp människor sätter på sig lager av kläder för den kalla vintern.
En kvinnlig bartender som serverar sina kunder ett leende, en dansare är i bakgrunden.
Kvinna bartender förbereda en drink med en pumpa på baren
En ung pojke försöker på underkläder som är för stora.
Två personer på en hockeyplan slåss.
En man med hjälm hoppar sin cykel nerför en trappa.
En man på en motorcykel omgiven av vit sand.
En grupp vandrare klungas samman på grå stenig terräng som gränsar till en glaciärs blåvita is.
En ung baseballspelare avrundar trea när utfältarna hämtar bollen vid staketet.
Unge pojke i en baseballuniform på väg att fånga en baseball i sin handske.
En man och kvinnor i orange på golvet skrubbning.
En publik tittar på två kvinnor klädda i traditionella asiatiska kläder förbereder sig för att skjuta pilar med sina bågar.
Fem män i hatt sitter i en cirkel och spelar olika horninstrument.
En liten pojke leker med en mopp som rör sig snabbt, och har många leksaker i bakgrunden.
En medelålders hockeyspelare som svänger på isen
En ung man rengör ett djur, medan två kvinnor ser på från bakgrunden.
En svart och vit hund som hoppar på en gård.
En basketspelare i vit uniform dribblar basketen mot en spelare i svart uniform.
Två kampsporter sparrar medan en domare med slips tittar på.
En kvinna som bär persikotopp och svarta jeans bowlar ensam.
Små indiska barn är samlade runt en bärbar dator.
En kvinna applicerar rött nagellack på naglarna.
En person bär svart skjorta och leker bowling.
En blondhårig flicka står framför en bowlingbana.
En ung kvinna målar ett tillkännagivande och ritar på ett fönster.
En ung man som hoppar från en brygga framför ett amerikanskt förortshem.
Hockeyspelare spelar ett spel på isen.
En löpare springer på en stig omgiven av gräs och träd.
En grupp åskådare ser Eiffeltornet från en balkong.
En man bowlar med olika nationella flaggor som visas i den motsatta änden på bowlinghallen.
Två äldre asiater som bär på en stor korg med produkter som de skördat.
Två pojkar på lek på ett roligt center, det finns två kvinnor i bakgrunden skrattar.
En man rider en wakeboard i havet.
Utföra några cykel underhåll, smörjer damen en ram innan monteringen är klar.
En man i blå skjorta fixar ett cykelhjul.
En asiatisk man i randig gul skjorta och shorts som bär lite kelp och vadar genom ett översvämmat område.
Ett rockband som spelar en livekonsert.
En person som bär hjälm och smutscykelutrustning rider en smutscykel över en kulle.
En dockteater som består av människor som står på höga käppar.
En liten blond pojke som bär en grön vinterjacka på stranden spännande tittar på vattnet.
En person som bär hatt sveper.
Två unga pojkar i badbyxor tvättar en stor brun hund.
En skridskoåkare snurrar på isen.
Pojken tar sin tur genom sprinklern och hoppar med glädje.
Cyklister rider tillsammans med trafiken på en stadsväg.
En kvinna som har tröja och keps chattar med en vårdgivare medan hon får intravenös medicin.
En man som bär grönt och svart hoppar genom luften och håller i en boll.
En bicyklist går sin cykel genom djup lera i ett lopp.
En liten afrikansk pojke ser nyfiken på en vuxen vit kvinna.
Två mörkhyade barn stirrar medan människorna bakom dem blandar damm i sina blommiga kläder.
En man i svartvit uniform spelar ishockey.
En man som bär headset spelar ett unikt instrument för en grupp åskådare.
En man och en kvinna lagar en måltid tillsammans i ett restaurangkök.
En svart man med grått hår, en vit skjorta och blå byxor sover.
Ett litet barn i gult och lila scooping småsten och smuts i en hink.
En fullsatt stadion vid 49-talets fotbollsmatch, med trupper som sprider ut en flagga.
Flera vuxna med gula hjälmar och flytvästar är forsränning.
En man med turkos väst och svarta byxor sätter sig framför ett tegelmonument.
Fem personer faller i skyn med fallskärmar.
Två afrikanska barn med ansikte målat i orange poserar för en bild framför en hydda.
En man i röd skjorta är bergsklättring.
En kvinna skalar ett svårt rockansikte med hjälp av ett rep.
Tjejen som spelar baseball bär blått och rött på ett basebollplan.
En ung hejaklacksledare uppträder med en trupp under en match.
En man i cowboyhatt sjunger och spelar gitarr.
En man som bär en mörkblå t-shirt och blå jeans och en yngre kvinna som bär en röd blommig klänning dansar tillsammans.
En man och en kvinna dansar medan folk tittar på.
En man och en kvinna som dansar ensam mitt i en folkmassa på en fest.
En ung kvinna åker skridskor på is.
Två kvinnliga skridskoåkare, en med mörkblå böjda uppåt och den andra med ljusblå böjda nedåt.
En barberare putsar en kunds mustasch.
En man som försöker slå sin golfboll som sitter fast i en sandfälla på en golfbana.
En individ hoppar över några jordramper på en svart och röd fyrhjuling.
En kvinna som bär en ljus, blommig klänning och en svart topp sitter på marken bredvid en byggnad.
En hane hoppar över vitt vatten.
En snowboardåkare flyger i luften och försöker landa på en snöhög.
En man i gula byxor är snowboard.
En blond kvinna i röd t-shirt och ett suddigt armband sjunger in i en mikrofon mot en grön bakgrund.
En person som hoppar högt i luften på en snowboard.
En motorcykelcyklist, klädd i full racingutrustning, kör över toppen av en sanddyn.
En manlig lärare undervisar sin klass av små barn.
Sex personer i tank toppar och hjälmar är rullskridskor medan två domare tittar på i bakgrunden.
En skidåkare är mitt uppe i att utföra ett mellanspel.
En ung flicka fotograferar utsikten nära skogsområden medan hon bär en sommarskjorta.
En byggnadsarbetare på en mekanisk lyft.
En ung pojke och en äldre man använder en övning på något slags föremål.
En ung pojkes färger på små pappersark.
En liten flicka som gör konst och hantverk med små paraplyer och korkar.
Barn gör hantverk vid ett hantverksbord med en vuxen.
Ett barn gör en aktivitet som involverar en cirkulär skiva med utstrålande linjer på den (i rött och blått, en limsticka, och utskurna nummer.
Ett litet barn lär sig om elektricitet med ledningar.
En elektronisk apparat håller på att arbetas på av en kvinna.
Ett barn interagerar med ett elektroniklaboratorium.
En man klamrar sig upp ur ett hål i isen upp för en trästege.
Två lag spelar hockey i en stadion, laget i gult gjorde bara en poäng.
Två hockeyspelare en i gult och en i vitt tävlar mot varandra för att få kontroll över hockey pucken.
Två spelare på ett fält slåss mot varandra.
En man som bär glasögon sitter i baksätet på en bil och spelar gitarr medan han tittar ut genom fönstret.
En man som hoppar för att göra en basketboll shot.
En grupp män spelar basket på en stål- och kedjebana.
En kille som åker skidor nerför ett berg i röd skiddräkt.
En college basketspelare stiger för ett hopp skott medan den motsatta spelaren försöker blockera skottet.
En motocross ryttare bär orange utrustning är turning ett hörn på kursen.
Två manliga hockeyspelare från motsatta lag är poserade på isbanan med sina hockeypinnar redo.
En ung kvinna hoppar sin häst i tävling nära havet.
Någon som bär gummihandskar tvättar disken i en metallsänka.
En kvinna uppträder med två hulahoops för en publik.
Folk tittar på föremål som visas på ett museum.
En pojke i röd skjorta leker med leksaksbåtar.
En person som bär en blå ryggsäck går upp för en snötäckt kulle.
Tre musiker som spelar för en sittande publik.
En man som bär en extremt kort slips, hängslen och färggranna randiga strumpor står på en scen och gör något med en anordning som involverar föremål som rullar fram och tillbaka på strängar.
En man med snöskor springer genom snön.
En hockey målvakt är på väg att fånga en puck.
Inga manliga byggnadsarbetare i ett arbetsområde i en stad.
Två barn, en bär blått, den andra bär rött, tävlar om att få en boll i ett spel.
High school basketspelare gör ett hopp skott med två spelare försvara korgen.
Två damer sitter på något som är gjort av betong, medan de njuter av ett mellanmål.
En tatuerad kvinna som klickar på en mus på ett skrivbord.
En liten flicka som poserar för kameran, uppklädd.
En kvinna i en park med ett rött paraply hoppar i luften.
En långhårig man tar ett foto av en strand.
2 personer, en i vitt, en i blått i en match
Basketspelare i orange uniform försöker blockera skottet på spelaren i den vita uniformen.
En gentleman i en vit labbrock kikar in i ett mikroskop.
Folk sitter på en strand och tittar på vattnet, med en man på en monter märkt Pipe Challenge.
Swans samlas runt en man och en båt.
Kvinna med glasögon, plasthandskar, och en labbrock, sätter droppar i ett provrör.
Ett barn dricker genom ett sugrör på sin dagis.
Kinesiska-amerikanska klädda barn klädda i röda uniformer gör en kulturell föreställning i en parad.
Två kvinnliga barn ligger i ett bad tillsammans.
Ett team av våldsamma hundar drar kraftigt en släde genom snöiga förhållanden.
En man skär deg i små fyrkantiga remsor.
En scen under ett hockeyspel där målvakten försöker hålla den andra spelaren från att göra poäng.
En man med glasögon som håller en nästan tom tallrik.
Två kvinnor spelar softball medan en bär lila glider till basen medan den andra bär vit försöker fånga en boll.
Studenter utövar yoga i en klassmiljö.
En man i en belamrad motorbåtsrad medan hans kvinnliga passagerare ser besviken ut i ansiktet.
En spansk kvinna bär en tung röd väska över axeln.
En grupp människor tränar på en gård och har händerna på huvudet.
En gitarrist framför musik på scenen.
Lilla pojke försöker hjälpa mamma att diska &amp; spela i bubblorna.
Två män, en som spelar horn och den andra som spelar sax på en svagt upplyst scen.
Två kvinnor klädda i röda zigenarkläder dansar runt i mörkret.
En blå tävlingsbil står parkerad på vägen.
Violinist spelar med bandet när det gula ljuset sätter stämningen.
En målarkonstnär pulvriserar en hona.
Man kan se två människor springa på stigar med träd mellan sig.
Denna rodeo idrottare försöker rida denna vilda häst.
Kvälls fotbollsmatch med ena sidan på väg att göra mål.
En ung man i röd skjorta får håret putsat.
Två personer trampar genom snön i ett terrängfordon.
Två killar i svarta jackor som använder och lyssnar på en skivspelare.
Flera män sitter medan de bankar på en bongo.
En liten pojke täcker sitt ansikte medan han är vänd mot lådorna.
Fyra killar i rullstol på en basketplan två försöker ta en basketboll i luften.
Två brandmän som slår på vattnet i slangarna.
En ryttare drar en wheelie på en motorcykel.
Två unga pojkar klädda i snödräkter leker i snön.
En man i blått med svart och gul väst spottar eld på en renässansmässa.
Två unga pojkar pratar med varandra.
En pojke med blå skjorta som leker på gatan med en leksak.
Isåkning ras går runt en kurva.
Tre vandrare vandrar i ett berg fyllt med träd och snö.
Fyra män springer på ett spår inuti.
Idrottsmän springer på en inomhusbana bär olika färgade skor.
Man på båt drar en lina från vattnet.
En tonåring i en blå Hollister märkeströja justerar ett "Sky-Waker" teleskop.
Surfare surfing i en vacker med fåglar runt och vågor med vacker textur
Ett lag av pojkar spelar basket i ett gym som en fan tittar på.
Tre spelare deltar i en lagsport.
En pojke med svart jacka och blå hatt kramar en brun och vit hund på en veranda i snön.
Byggarbetare arbetar på en scen.
Fyra clowner, två män och två kvinnor, går nerför gatan och vinkar.
En pojke hoppar en cementvägg med en grön skateboard.
En man rider en orange skateboard i en skateboardpark.
Lilla flicka som leker klä upp sig i rummet bredvid sina leksaker.
Turisten använder kikaren för att få en bättre utsikt över det fridfulla havet.
Spelarna är i sin dagliga rutin träning.
En dykare ignorerar en grupp blå och gula fiskar när han utforskar havet.
Tre dykare kommunicerar med varandra.
En man i grön skjorta, stående på en kanna hög har precis kastat en boll.
En kille undersöker något under ett mikroskop medan folk tittar på.
En hane i blå jeans och en blå skjorta som jobbar på några inomhusstolar.
Fem arbetare i orangea kläder och blå hjälmar arbetar med byggnadsställningar.
Man i vit karate uniform, vänder en annan person i en blå uniform med folk som tittar på.
Två pojkar i brottningsmatch.
En asiatisk ungdom som sitter på en vägg med en skateboard i knät.
En stråkkvartett busking för en publik på gatan.
En man i svart läderjacka spelar saxofon.
Ett barn står upp och ner i en pool.
En liten flicka borstar tänderna framför en spegel i badrummet.
En man som håller i en gitarr sjunger.
En man jonglerar flammande föremål med ett staket och en bil i bakgrunden.
En liten hund som leker bogserbåt med en större hund
Över huvudet på två personer, en man och en kvinna, som tillagar en måltid med potatis.
En man i grå skjorta som spelar fiol.
Ett barn i grön jacka rullar en bowlingboll mot stiften i sin fil.
En liten pojke som bär en Marvelskjorta borstar tänderna.
En äldre man cyklar med en blå tvättkorg full av kläder på styret.
En kvinnlig skidåkare i en blå tröja ler ovanpå en stor kulle.
En man som bär en stor ryggsäck navigerar sig fram genom snötäckt terräng.
Två killar som monterar en låda på ett räcke.
Ett lag av Roller Derby Girls blockerar tävlingen när de går för segern.
En man klädd i snödräkt åker längdskidor.
Unga manliga soldater i kamouflagebyxor och hjälmar städar upp skräp utanför en byggnad.
En hockeyspelare i uniform sitter på en hockeybana.
En skjortlös man med en kapplöpningsskylt på rumpan poserar som en kroppsbyggare.
En pojke hoppar 5 trappor på en hopfällbar scooter.
Damen med en vit handduk på huvudet säljer på en öppen marknad.
En grupp unga män klädda i rött går förbi en turnébuss.
En man i jeans och en knapp upp skjorta presenterar något på en projektor skärm.
Två män är på en båt och tvättar vattnet.
En bartender med vit skjorta häller upp ett glas apelsinlut.
Person klädd i tidningspojkkläder som häller upp drinkar.
En man i randig skjorta, väst, slips och hatt serverar sig själv slag från en stor skål.
Någon släpper orange mat färg i en klar drink.
En bartender med en svart knapp upp skjorta häller två drycker.
En bartender skakar om en drink.
Två män, en i svart och en i grått, utför ett vetenskapligt experiment.
En kvinna som blandar drinkar i en bar och poserar för kameran.
Tre personer, två män och en kvinna, poserar för en bild med flaskor med drycker och klädda i vetenskapsklänningar.
En äldre man och kvinna är redo att manövrera en apparat.
En kvinna som besöker någon form av konferens skapar ett projekt på en iPad.
En man i rutig skjorta säljer produkter till kunderna.
Man i vitt och rött tackling man i grön skjorta för bollen.
Folk är redo att ta en gul buss.
Tre personer på motorcyklar rider ner på en grusväg.
Två surfare, en skjortlös, rider en våg.
En flicka med svart vinterjacka och bruna stövlar kastar snö över ett staket runt en kanal eller vattenväg.
En man i hatt och overall förbereder en god maträtt.
En man på en trottoar i en rock som spelar mässing klarinett.
Tre vänner dricker kaffe.
Det sitter folk på en buss och kameran är fokuserad på en man som viftar med händerna mot kameran.
En grupp människor klädda i badkläder står utanför i ett snöigt, skogsaktigt läge.
2 hockeyspelare i svart guld och vitt, en har pucken med sin pinne och är skridskoåkning.
Fyra damhockeyspelare rusa efter en lös puck när det hoppar längs brädorna.
En person på en smutsig fyrhjuling som kör genom jorden.
En skjortlös äldre man som gör en traditionell indisk gatumaträtt.
En man i röd skjorta ger ett fredstecken medan han lagar kyckling på en grill.
En man och en kvinna som tittar på ett barn.
En ung man ligger under ett stort träd i en park och håller i vad som verkar vara en öl.
Brandmän står på taket av en byggnad omgiven av träd.
Två män i uniform drar i en stor kabeltråd.
En man i mitten av ett hopp medan snowboard.
En snowboardåkare slipar på en skena nerför en sluttning med snö runt omkring.
Tre herrar spelar basket, en man med bollen och två försvarare på sig.
Två små barn i svarta kläder och stoppning utför en kampsport match där de tävlar mot den andra.
En rad gamla vagnar dras av boskap.
Du afroamerikanska pojke utan skjorta på leende medan hålla en skål med mat.
En mountain bikeer är i luften mitt i ett stunt.
11 män och kvinnor sitta runt ett bord äta, medan 1 kvinna böjer sig över i bakgrunden.
En kvinna med röd halsduk jonglerar med apelsiner.
Ett lag är hopblandat på spelplanen, bär blå skjortor och blå och röda shorts.
En man i ljusa färger får hjälp att utföra sina rutiner.
En fotbollsspelare bär en röd och vit uniform fånga bollen för en poäng som motståndaren bär en blå och vit uniform är i bakgrunden tillsammans med en mängd människor tittar på spelet
Flera fotbollsspelare i defensiv position (s ) på marken under ett spel.
En man i blå byxor står bakom en bil parkerad på gräs utanför en tegelport.
Ett barn i tröja och jeans kjol hukar.
Fotografen fångar sin skugga när han fotograferar unga pojkar som minglar på gräsmattan.
Folk i parken tittar på matchen.
Den här bilden är av en man i en udda dräkt som jonglerar.
Två personer är utanför och grillar lite kött.
En person på en skidbräda tycks ha hoppat från den närliggande helikoptern.
En man som hoppar på en skidbräda.
En man spelar ett instrument på en konsert.
Ett par kvinnor som bär tegelstenar på huvudet.
En person i solbränna och blå tröja hängande kläder på en klädstreck utanför fönstret i hennes byggnad.
En kvinna mitt i kastet av en bowlingboll.
En grupp små barn skrattar och leker mitt i stora bubblor.
Kvinnan pratar med en fotograf klädd i svart.
En skäggig man i solbränd hatt, hjälper en skallig man i tennisskor, nära en lägereld.
En kaukasisk hane i en grön och vit rutig skjorta som håller en mikrofon.
Män och kvinnor med väskor och portföljer reser upp och ner svagt upplysta rulltrappor.
Fyra inomhuscyklister tävlar runt en krök.
Fyra cyklister, tre av de in-line och en till sidan, cyklar längs banan.
Basketlag, med en av spelarna på väg att gå för ett skott.
En grupp unga män som spelar basket; två medlemmar i samma lag försöker blockera en spelare i det andra laget som har bollen.
En röd och vit bil rundar ett hörn på en kapplöpningsbana.
En person som går i snön med en skog av träd i bakgrunden.
En kvinna skriker in i en mikrofon medan hon bär en röd jacka.
Två spelare möter ishockey som domaren har just kastat pucken på isen.
Två män i röda skjortor och blå byxor spelar hockey.
Två svarta hundar slåss framför en solbränd soffa.
Jag har verkligen ont efter att bollen studsade från pannan.
En kvinna som bär en bricka med drinkar på.
En kvinna är helt täckt och fixar en maskin.
En man med en gul hård hatt på arbetar över lite vatten.
En kvinna som sitter i hörnet och bär en blå rutig sjal.
En kvinna ligger i sängen med sin katt när hon husdjur henne.
En man förbereder sig för golf, och det finns en stor publik som tittar på honom.
En man som tittar på någon form av contraption medan en annan man i bakgrunden tittar på.
Kvinnor som visar ett barn hur man löder en metallbit.
Två små barn använder en mortel och mortel slipning en produkt ner.
En kvinna visar ett barn hur man använder en symaskin.
En ung flicka i rosa skjorta skapar en målning på papper.
En ung man i blått som arbetar med elektronik.
En man maler en bit metall framför en åskådare på en studio.
Protestörer håller skyltar på spanska.
Två män, en med mohawk och solglasögon kryper genom leran, medan andra ser på.
En musiker klädd i kostym spelar sitt stora instrument medan han sitter på en förstärkare.
En pojke i blå skjorta är på en skateboard i luften gör stunt, medan andra tittar.
En cykelförare med en kostym täckt i annons förbereder sig för ett lopp.
Flera män i gul och grön väst i ett café som äter lunch.
Två basketspelare i vit tröja vaktar en spelare från det andra laget.
En person med glasögon och en svart mössa böjer sig över utrustning i mörkret.
En snowboardåkare tar flyget medan han utför en fristilsrörelse.
En blå-röd och huva figur går förbi ockuperade bord i ett överklass rum.
Detta en man på en båt i lugnt vatten omgiven av träd.
En liten flicka står på trottoaren och blåser bubblor.
En man utanför Rodgers slaktare tittar på mat.
En man lutar sig mot en eld för att kontrollera innehållet i en gryta.
Soldaten hoppar från planet
Två unga flickor i klänningar hula hänger på gatan.
Stenar utanför sitter i solljuset och kyler sig när solen går upp.
Män leker med en volleyboll i en pool.
Tröjlös man som spelar tangentbord och sjunger in i en mikrofon.
En leende kvinna och fyra små barn som poserar för en bild.
En man och en kvinna poserar tillsammans framför en vattenförekomst.
Två unga flickor kysser en man på vardera sidan av hans ansikte med en fyr på en kulle som bakgrund.
En pojke och en flicka ler för ett foto medans de är i en pool.
En snowboardåkare som sparkar upp snö under ett träd på ett berg.
En liten pojke i blått har ett gult föremål framför en blommigt designad stol.
Ett rugbylag jagar när mannen i besittning puntar bollen.
Män spelar hockey på rullskridskor.
En asiatisk frisör med en handduk över armen står bakom en tom frisörstol.
Två män med ansiktshår som gör tortillas i en informell miljö.
Ett postbolag med ett stort leende står på trottoaren med sin postvagn.
Mannen blir kysst av två vackra kvinnor.
Två tonårspojkar övar sina fotbollskunskaper när deras vänner står bredvid målet och tittar.
En kvinna i en blå klänning står med en skamlig min i ansiktet.
En man med grått skägg i karateläge med ett gult bälte på midjan.
En liten pojke i röd hatt med en Ritz kex i handen.
En kvinna i vit blus skrattar, medan en annan kvinna i svart skjorta och glasögon ser på.
En kvinna ler när hon ger en presentation på en mikrofon.
En ung vit pojke som står ensam i ett rum och jonglerar med oidentifierat material.
En man i uniform hälsar.
En man spräcklig med blå, orange och grön färg över sin överkropp håller upp en kamera.
Människan skyfflar smuts i en hög
Människor från alla samhällsskikt rusar för att hinna med nästa tåg i Japan.
Små barn leker med hulahoops i ett stort rum.
En kvinna i ett svagt upplyst rum tittar genom sitt mikroskop och justerar synen.
En löpare deltar i en löpning eller tävling längs en ödslig sträcka av landvägen.
En familj väntar bredvid några bärbara toaletter i staden.
Två killar som jobbar utanför räcket.
En man i en olivgrön skjorta som använder en hammare för att skulptera ett gyllene föremål.
En familj på fyra sitter på ett täcke i en skara andra.
Flera personer med ljus runt omkring eller i handen är vända mot kameran eftersom de var och en har olika antal fingrar som hålls upp.
En man jonglerar tennisbollar bredvid sina två vänner.
En vit man i ett vitt rum fylld med bilder som sitter ner och försöker sätta ihop en ram.
En säljare som bär ett rött förkläde och säljer mat på en fotbollsmatch.
En basketspelare i en gul uniform försöker dribbla medan han försvaras av en spelare i en blå uniform.
En flicka skrattar medan hon sitter på en soffa.
En man hjälper en liten pojke att klättra upp för en stolpe som finns på lekplatsutrustning.
En svart hund som springer mot kameran.
En ung man spränger vattnet i ett par glasögon i ansiktet.
Två unga män i uniform deltar i en basketmatch.
En kvinna sveper utanför ingången till en byggnad med två stora trädörrar.
Två spelare möter i en basketmatch.
En kvinna som bär solglasögon, en röd skjorta och svarta shorts springer i en road race.
En mans huvud blir senare efter att ha klippt sig.
En man med glasögon och rött ansiktshår berättar en historia för två leende män.
En man med skägg håller ett par tångar vid ett restaurangbord.
En man med skägg och overall står bredvid två män med svarta jackor.
Ett barn med blå ögon och ett smutsigt ansikte pekar på hans vänstra öga.
En äldre man som bär skridskor och håller i en hockeypinne tittar på en hockeypuck i luften.
Den här unga flickan tar sig hem.
Det finns människor på en golfbana och en dam håller en flagga vid ett av hålen.
En liten pojke i hatt som plockar upp påskägg.
Två män med motorcykelhjälmar, en med papper.
En blå hiss som sätter upp dekorationer på en byggnad.
En man surfar och är i luften med vågen plaska bakom sig.
Två personer som bär hjälm cyklar i skogen.
En man med vit hatt och verktygsbälte som jobbar på taket.
Två män med hattar som spelar ultimat Frisbee.
Två killar, en i vitt och den andra i rött hoppar för att fånga en frisbee.
En man gör en dykning fångst under ett spel av ultimata frisbee.
En man i vit t-shirt och khakis har en fantastisk eld jonglering show.
En mager pojke flockas i smutsigt vatten med sina smala byxor.
En vit och gråfärgad häst hoppar ett gult tävlingsstängsel medan dess ryttare håller i sig.
Två poliser patrullerar på sina hästar.
Ett fotbollslag är på en spelplan, några av dem fixar näten och en tömmer vatten från en kylare.
Medlemmar i ett fotbollslag kramas på fältet.
Fotbollsspelare är på ett fält, en på väg att sparka en boll, och en annan försöker stjäla den från honom.
Fyra fotbollsspelare tittar på en boll, två styck på separata lag, som nummer 10 Messi sparkar bort den.
Ledaren var mycket upprörd under föreställningen.
Tre personer är synliga deltar i sporten fäktning medan två åskådare tittar bakifrån.
Det finns ett team av vinteridrottare som skidåkning tillsammans i en linjeformation.
En person som tvättar händerna i ett vitt handfat.
En Roosevelt fotbollsspelare röv huvuden med bollen och en motståndare under en match.
En hastighetscyklist går runt ett spår med domare som observerar.
En man som bär cowboyhatt, overall och vit skjorta pekar på sitt musikark och tittar på någon som är förvirrad.
En rallybil driver runt en sväng och stänker lera.
Tre vuxna, två män och en kvinna som pratade med varandra på vintern i snön.
En grupp ungdomar klädda i uniform går nerför gatan.
Ett barn i gult försöker ett mål på en fotbollsmatch medan målvakten i rött försöker blockera skottet.
Gentleman gör en pjäs på en fotbollsboll
En pojke i gul huvtröja och en flicka i rosa kläder leker på stranden.
En vit man undervisar en klass i Asien.
En blondhårig bebis klädd i rosa och vitt håller i en tandborste.
Flera svarta barn är samlade poserar för bilden i ett fält.
Blond kvinna i rosa skjorta borstar en brun häst med vagn hjul i bakgrunden.
Det finns en liten flicka i en rosa skjorta som håller en röd handväska i handen
En person krossar ett ägg i en silverskål med bara en hand.
En baseballspelare glider in i andra basen medan motståndarna hoppar infielder.
En man som står längst fram i rummet pekar upp medan flera människor som sitter tittar mot honom.
En manlig publik på en strand kastar sig bakåt när man knäböjer i mitten.
En hund är avståndet hoppa i en pool av vatten medan åskådare tittar.
En man i svart skjorta blandar drinkar
En man skateboard på en bänk bredvid ett böjt träd framför en vit byggnad.
En man och en kvinna är ute på fältet och håller varandra i handen.
En grupp barn står vid ett barnbord och stolar medan en av dem sätter sin fot i en liten plastbehållare.
En brun hund springer genom fältet.
En basketspelare i en St Johns nummer 10 jersey doppa en basketboll.
En skidåkare i röd sprayar snö mot vit bakgrund.
Dessa kvinnor njuter av det fina varma sommarvädret i det tropiska samtidigt som de njuter av en uppfriskande drink.
En man i mörk jacka jobbar i en träaffär.
En äldre kvinna försöker på en svart hatt medan hon tittar i en spegel på en klädbutik, med en försäljningsassistent till höger.
En djärv motorcyklist som zoomar genom en kapplöpningsbana.
En kvinna ritar vid ett bord med en blå permanent markering.
En ung flicka med en handritad klocka pratar med två kvinnor.
Liten asiatisk flicka med gula glasögon arbetar på en bit träarbete med hjälp av en vuxen.
Baseballspelare och umpire på hemmaplan gör en pjäs.
En man med lila mönstrad skjorta och jeans sitter på en brun rekyl.
Två motorcyklister tävlar på en asfaltbana på lila och gröna motorcyklar.
En grupp tittar på en man i vita byxor med en yxa.
Två go-cart förare tävlar på racerbanan.
En person på en cykel hoppar över gräs och stenar på en utvändig stig med ett berg i bakgrunden.
Två män spelar fotboll på ett plan.
En hand syns hålla en liten sil med en röd substans inuti.
Kvinnan njuter av att ha en annan beskyddare bakom sig.
En man håller sig i nosen medan han smakar på något och kvinnan skrattar åt honom.
Grupp av barn och en vuxen man som ligger på golvet med bollar på huvudet.
En kvinna i bikini och solglasögon stöter på en volleyboll på stranden.
Blake Griffin, av Los Angles Clippers dunkande över en Minnesota Grizzles spelare.
En man klädd i svarta byxor, en orange och brun randig skjorta, och en svart bandanna i en "bara kastat en bowlingboll" ställning.
Ett band som sjunger för en massa människor.
En grupp män och kvinnor arbetar på olika delar av viktlyftningsutrustning.
En man sitter bakom ratten i en bil.
En ung pojke, klädd i cowboykläder, rider en galopperande häst.
Manlig idrottare i luften, bär vita shorts och höga topp skor.
En Marquette University spelare går mot korgen, och ifrågasätts av en St Johns försvarare på Madison Square Garden under Big East Tournament.
En man drar i en kedja i en verkstad.
En ung pojke i grå hatt, klädd i mestadels svart, tar emot skosnören och spelar på skateboarden.
Två unga, manliga fotbollsspelare tävlar om bollen på ett vått fält.
En tjur försöker kasta av sig en manlig människa med färgglada byxor på ryggen.
En man, i röd skjorta, rider på en gammal traktor.
Ett litet barn i en röd jacka som rider på en kvast som en häst.
En man och en kvinna klädd i vitt övar elddans.
En musiker i en enkel grå tee knäböjer framför sina trummor på en plankscen i trä.
Mannen bär en ljusblå jeansjacka och tittar på en målning bredvid en flod och bro.
Lilla blonda tjejen i jackan sticker ut tungan medan hon håller i en röd ballong.
En hund i gräset framför en byggnad.
Två kvinnor på rullskridskor med hjälmar och armbåge och knäskydd stöter varandra när de skakar.
En spektakulär dunk av en professionell spelare med vit och gul på
En svart man i vit uniform gör en spektakulär omvänd smäll till publikens förvåning.
Ett asiatiskt par som bär blå och röda formella kläder står tillsammans i en skogsmiljö.
Två män bär vita kläder och hjälmar är forsränning i vitvatten forsar.
Skidåkare och snowboardåkare värmer sig vid elden medan de pratar.
En depå besättning reparerar till en motocross cykel medan deppbesättning chefen övervakar.
En kvinna som sitter vid vattnet och tvättar lite kläder.
En pojke gör en vända medan en annan pojke står på Matt.
En kvinna läser bredvid en vattenfontän.
Tre damer nära ett bord utspridda med böcker, upptagna med att skriva anteckningar från sina referensböcker.
Tre tjejer som spelar hopprep utanför.
Två män sitter på ett café och pratar, medan en suddig kvinna i en lila ytterrock går förbi.
Två afroamerikanska män tränar på en fotbollsplan.
En man sitter ute i den partiella skuggan i en hängmatta och läser något.
Två män för ett samtal på en trottoar.
En ung man försöker sticka valv över en bar, knappt några centimeter bort från den mitt i flygningen.
Den här hunden verkar inte uppskatta hur grym hans hatt är.
Hunden sitter på soffan med ett julband ovanpå huvudet.
En kvinna med ett riktigt smutsigt kök som diskar.
En kvinna med kort hår i kjol, skjorta och solglasögon jonglerar med tre apelsiner.
En man som strör majsen på marken.
En spelare från Oakland A: s glidande till andra som spelare från Änglarna väntar bollen.
En basketspelare avvisar en annan basketspelare skjuten i luften precis under korgen.
Två branta hästar, kör parallellt, gör ett hinder språng, på banan med sina ryttare.
Det är en vacker dag på hästkapplöpningen.
Två jockeys leder sina hästar över ett hinder under ett lopp.
Bröd delas mellan en man och två kvinnor.
En man som håller upp ett ljust rosa paraply på en stadsgata.
En kvinna arbetar som sömmerska.
Kul kille leker med sin mjölk halm ger ett leende för kameran.
En motorcykel racer tar en tumla medan två konkurrenter kommer racing upp snabbt bakifrån.
En snowboardåkare utför ett trick genom att rida nerför rälsen i en trappa.
En liten pojke leker med en skateboard.
Fotbollsspelare i vitt och grönt dyker för bollen som han försvarar mot sin motståndare i svart.
Hockeyspelare tar pucken.
Ett lag av män spelar ett spel där flera av dem hoppar för att nå bollen.
En man tittar på en gul bulldozer.
En bulldozer skjuter stenar och smuts i en hög.
En gul bulldozer maskin i ett stenigt fält.
En gråskäggig man skär blad i några fjäderfän på en skärbräda.
Unga flickor samlades runt en man som blåste stora bubblor.
Blå och grå segelbåt i vattnet med några andra båtar framför mot en grå himmel.
I det här fotot har vi två fotbollsspelare som går för en rubrik.
En man som ligger ute i skuggan av ett träd med solglasögon på medan han läser en bok.
En man kollar sin telefon medan han sitter på en stenbänk.
En skara människor som ser på som en stor staty av en man flyttas.
En man fångar en stor våg på sin surfbräda.
En tjur sliter av en ryttare som bär en rosa skjorta och chaps.
Ett litet barn i en baby sving som har en gul klänning på sig.
En Atlanta baseballspelare bär en handske på infältet.
En ny pappa ser att hans faderskap fortsätter.
En man på en mountainbike rullar nerför en mild kulle.
O Åh cool gå gyttja, fick min hjälm och jacka.
Ett litet, blont barn klappar en liten hund utanför.
En ung gymnast övar innan en match.
En ung man i blå jeans och en blå tee-shirt en solglasögon är på en skateboard på trottoaren kantad av palmer.
En kvinnlig sångare och manlig gitarrist och trummis uppträder på en scen.
En kille med öronmuffar och skyttar glasögon placerar gevärets sikt på ett mål.
En man som övar på att skjuta med sin säkerhetsutrustning på.
Tre shortboardare går nerför stranden mot en våg av svarta stenblock.
En man står i kokosnötter och försöker öppna en.
Många människor av alla raser är samlade omgivna av röda, vita och svarta ballonger.
En kille i sin dykutrustning pratar med andra män.
En grupp barn som spelar fotboll av ett gammalt slott.
Det finns en grupp människor på en traktor av något slag som rider genom ett fält.
En man, i en svart kortärmad logotypskjorta, sitter vid en elektronisk konsol med hörlurarna på.
Kvinnan bär en blå tröja samtidigt som hon håller i en stor bit brunt pappersmaterial.
En kaukasisk kvinna med blont hår och en rosa rosett lägger ett föremål i en plastpåse.
En man som cyklar genom lera i full kostym.
En man med blå hatt och svart väst rider en brunfärgad tjur som sparkar upp damm.
En skidåkare hoppar en snödriva högt i träden.
Gör allt klart för publiken på den spanska matrestaurangen i NY.
Ett team av tjejer som tävlar på rullskridskor.
En man klädd i en surfskjorta och blå och vita shorts guidar skickligt sin gula bräda med dess mångfärgade segel över krönet av en havsvåg, vänder sig över i processen.
En basebollspelare har just slagit bollen och är på väg att springa.
En fotbollsspelare i en grön jersey sparkar en blå och gul boll.
En liten pojke i hjälm och klädd i svart, svänger en blå fladdermus i tee boll.
En kvinna som tar en bild medan hon njuter av ett glas vin.
Tennisspelare återvänder en hög serve på tennisbana.
En man verkar sy något slags material.
Fotbollsspelare i sina uniformer kör upp fältet mitt i ett spel.
En pojke med armen inlindad i ett ACE-bandage vilar i en säng.
En ung pojke är mitt uppe i en försäljning av getter
En man och en kvinna i jeans sitter på båda sidor av en gitarr.
Två brottare brottas i ett gym.
En hockeymatch pågår i en stor ishall.
En man regisserar en kamel som bär på lite material.
En konst- och hantverksklass målar ett projekt medan läraren övervakar och ler mot dem.
En man i en basketmatch skjuter bollen.
En grupp unga människor sitter runt en brandgrop.
Tre spanare är på toppen av en klippa med utsikt över havet.
En man försöker sätta dit sin motståndare som krigar mot en blå singel under en brottningsmatch.
En man i hjälm och uniform ler.
Många cyklister är redo för en tävling.
En man som har ansiktet täckt med en turban bär ett vapen.
Glidande nerför en snötäckt kulle på en släde, med träd och berg i bakgrunden.
En liten flicka med ett stort tecken som säger "END WAR" och hon tittar ner på det.
En tabell full av gymnasieungdomar utför vetenskapliga experiment i tre grupper om fyra.
Studenter undersöker foton på nära håll i klassen.
En pojke rider en leksakshäst, som placeras i hörnet av en teal tegelhörna.
Arbeta med att borra på trä för att göra hål.
En målvakt spelar hockey, och det finns ett objekt framför nätet.
Fem personer sitter runt ett soffbord och går igenom lite pappersarbete.
En svart hund springer på grönt gräs mot kameran.
En skallig man är på en surfbräda antagligen redo att fånga några vågor.
En man i sitt kök lagar en god måltid.
En manlig sångare spelar gitarr och sjunger under strålkastarljuset.
Tre personer klättrar i matchande kläder bredvid ett litet vattenfall.
En man spelar trummor.
En mörkhårig man surfar från en stor havsvåg och är luftburen.
En man på en atv njuter av en eftermiddag ridning i öknen
Tre personer står stolt vid en lastbil fylld med byggnadsmateriel på gatan.
En man i goggle som simmar.
Ryttare i rött racing en mini röd racerbil som rider mycket nära marken.
Två barn och en vuxen som gräver ett hål i sanden i vinterkläder.
En asiatisk kvinna, klädd i en ljusrosa skjorta, tvättar sina kläder i floden.
Snöskidare flyger högt genom luften.
En person i orange byxor åker skidor nerför en sluttning.
Två tjejer som leker inne i ett hopphus.
En djuphavsdykare är i full utrustning och studerar en havssköldpadda.
En man med en gammal kostym som dansar i en balsal med en kvinna.
En kvinna i en ljusrosa kjol som bär en korg på ryggen och går uppför en kullerstensstig.
En person som går längs en väg i öknen.
En man har just vunnit från en karatestrid med sin motståndare och hans näsa blöder.
En äldre man, klädd i salongsdraperi, klippt sig.
En kvinna med en röd luva som försöker korsa en ström av vatten skolös med en täckt TV.
En flicka med leopard knä hukar medan rullskridskor nerför banan.
En manlig hejaklacksledare håller en kvinnlig hejaklacksledare i luften på en fotbollsmatch.
Människor med anti-immigrationstecken.
Ett litet barn, som bär randig skjorta, kan inte se nerför teleskopets rör.
En frisör klipper en äldre man utomhus.
Ett par män sitter utanför medan den ena spelar dragspel och den andra spelar ett vindinstrument.
En grupp människor hänger utanför.
Tre unga pojkar leker i sanden längs stranden.
En grupp indianpojkar som gav fredstecken.
Ett par går igenom öknarna i ett rum fullt av människor som är intresserade av mat.
En kvinna sitter på en soffa med fötterna uppstoppade på ett bord, medan hon använder en laptop.
Mannen försöker göra en keramik som han kan sälja snart.
Två indiska damer fotograferar det långa gröna gräset utomhus i sitt hemland.
En kvinna som får en ryggmassage från en man medan hon sitter på en basketplan.
En man och en kvinna utför kampsport utomhus.
En man som gör ett trick på sin BMX cykel på toppen av en halv pipa
Två män i en stad som arbetar på en byggarbetsplats, med höga byggnader bakom sig.
Det finns fem jockeys på hästar med träd i bakgrunden.
Två hockeyspelare står med båda armarna upplyfta.
En afroamerikansk man springer nära vattnet utan tröja.
Två män och en kvinna springer tillsammans för en tävling.
En skjortlös svart man som bär solglasögon och joggingbyxor längs en parkstig nära en vattenväg.
En arbetare som tar ett glas vatten.
Två män i blå uniformer och hattar tillsammans med vita stövlar går längs en gata.
Dessa män marscherar band spelar instrument på gatorna.
En kvinna på en restaurang lagar mat på en grill.
Reporter tar en intervju från en röd racerbilsförare.
1 killar springer med en vit boll fotboll i sand medan en annan jagar honom.
Fem militärer står framför en staty.
En man i en blå och orange skjorta sparkar en fotboll till sin lagkamrat.
En manlig idrottare slår huvudet i marken för att skydda bollen i lek.
På en urban marknadsplats får en man klippa sig med flera andra män och en liten flicka i bakgrunden.
Två killar lastar lådor i en blå behållare som sitter på en tegelpläterad gata.
En man gör en lerkruka, medan flera åskådare tittar på.
En man sparkar en boll på ett fält.
En man visar tre kvinnor hur man skapar keramik i en klass.
Den här killen har precis skapat ett nytt sätt att laga mat till sin familj.
Mäns Volleyboll lagets medlem hoppar upp i luften för att spetsa bollen i de andra lag som spelar planen.
En grupp kvinnor som lämnar ett hinder i ett lopp.
En man lägger sin första fot i en låda fylld med vatten.
En publik tittar på när sex män förbereder sig för att springa ett lopp.
En man med svart skjorta, röd slips och röda hängslen koncentrerar sig på att jonglera tre röda bollar.
Två killar som spelar fotboll på planen.
En ung flicka i leopardtryck står i köket och håller en spatel medan hon lagar pannkakor.
En man på en vacker strand använder en kniv för att öppna en kokosnöt.
En snowboardåkare tappar balansen och dyker ner i snön först.
Två män i blå skjortor som ler och skakar hand.
En kvinna i lila skjorta som springer ett maraton och får vatten stänkt på henne.
Många poliser i upploppskläder omger en man i vit skjorta.
En grupp ungdomar dansar med entusiasm med sina partners.
Flera människor väntar utanför på evenemanget.
Två idrottare, en med lila och blå ränder och den andra med blå och vita ränder, spelar fotboll på ett plan.
Man i gul skjorta utför underhåll på Schwinn cykel nära ett picknickbord.
En ung pojke bowlar för en nål med en boll utanför, medan tre andra personer är i bakgrunden.
En kvinna i en rutig kappa som äter sockervadd.
En företagspresentation där presentatören bär randig skjorta och använder en projektor.
Kaukasisk man i en hård hatt håller en kraftborr framför den amerikanska flaggan.
Barnet i en blå jeanshatt och solglasögon tittar på kameran medan det hålls.
En skäggig man i svart står tvärs över gatan från en Bradford's.
En rugbyspelare passerar bollen när han närmar sig en försvarare.
En grupp fiskare som håller ett nät och tittar på ett litet parti fångad fisk.
Flera män spelar hockey med åskådare sitter på läktare.
En arbetare städar ett tak eller en terrass på en kall vintermorgon.
Lödare i en marschparad som står stilla vid uppmärksamheten.
Två män utomlands tycker om att tala om sina olikheter.
En man med sin hund bär vandringsredskap och tittar på utsikten över bergen.
2 hockeylag spelar hockey.
En man i rosa skjorta står bredvid två yngre män i ett mörkt rum.
En liten bild som används för att beteckna en trasig webbbildlänk
En fotbollsspelare för Eik hoppar högt i luften för att sparka bollen, jagas av flera motståndare och en lagkamrat.
En kvinna som tittar på när två barn leker vid en pool.
Fyra kajakpaddlare i två färgglada kajaker "surfar" en stående våg i en flod som flyter genom en park.
En kvinna med svart klänning och solglasögon jonglera citroner utomhus.
En kvinna ritar en hund med blyertspenna på ett litet torg.
Ungt barn använder verktyg på en maskin.
Äldre man pratar med en ung pojke som bär en blå och brun skjorta.
En ung pojke förbereder ett projekt med en skäggig man.
En grupp på åtta personer som spelar någon form av bordsspel runt ett bord.
En ung flicka lär sig hur elektriska kretsar fungerar.
Barnen befinner sig i en klassrumsmiljö och lär sig att sy på en symaskin.
En person som väljer ett lås med en bit metall.
En ung flicka som bär färgglada kläder använder henna för att rita en blomma på handen.
En ung pojke i glasögon använder en hammare på ett metalliskt föremål.
En flicka visar upp vad jag antar är konst hon gjort.
En ung människa som tar isär eller sätter ihop en elektronisk apparat.
En ung pojke i en blå jacka tittar på något som sågas isär medan han bär skyddsglasögon.
Elementärskolans elever tittar på ett experiment i en stor glasapparat.
En man fångar en boll mitt i någon slags sport.
Tre personer springer genom leran med folk i bakgrunden.
En man i bruna kläder och sandaler sopar ett stengolv.
En äldre person öppnar ett glas och väljer en ost.
En basketspelare dunkar basketen under ett spel som publiken och spelarna tittar på.
Spring, spring försiktigt, slå inte på skåpbilen.
Två studenter på jobbet i en naturvetenskaplig klass.
Två flickor sätter en kemikalie i en flaska.
En brunett äter nudelsoppa med ätpinnar ur en orange skål
En person står på en stege och sätter upp bokstäver på en skylt vid en teater.
Ett stort vitt växthus med en familj som sitter framför det och har picknick.
Svart hövding gör en mat på hotellet
Fans och spelare firar och lyfter sin tränare på sina axlar efter att ha vunnit en fotbollsmatch under en nattmatch.
Två sexiga kvinnor brottas i ringen.
Vit man som spelar gitarr live på scen i ett rockband.
En ung flicka i rosa och zebra-tryck ler medan hon håller ett uppstoppat djur på en födelsedagsfest.
Ett barn i röd rock tittar genom linsen i ett metalliskt blått teleskop.
En ensam clown lägger till en välbehövlig färg till världen.
En vattenskidåkare dras av ett rep och han bär rosa och svarta byxor.
Två unga män inspekterar ett kar och rör på en hamn.
En mörkhyad man i vit uniform avleder en boll från målnätet.
En fotbollsmatch mellan ett lag med vita tröjor och ett lag med gula tröjor.
Fyra motocross racers flyger över off-road dirt ramp under en tävling.
En flicka i vit jacka ler medan hon håller i en mikrofon.
Fem ishockeyspelare från samma lag firar på rinken.
Män som spelar ishockey och en har just fallit.
En scen från ett hockeyspel där spelaren i blått just har tagit ett skott, medan spelaren i vitt försöker blockera det.
En pojke som håller en stor sten med en annan pojke suddig i bakgrunden.
Två barn, en flicka och en pojke, tävlar i ett potatissäcklopp.
Amish killen spelar golf och promenader
En kvinna i ett rött förkläde ser på när en man i ett svart förkläde knäcker ägg.
En kock på en enhjuling jonglerar genom en skara åskådare.
Det finns en flicka med tre pojkar som simmar i vatten.
Kvinnlig distanslöpare deltar i ett lopp.
Fem män, klädda i orangea reflekterande kostymer, arbetar på järnvägar.
En man med glasögon som jonglerar för barn.
En baseball man glider sig till basen medan den andra mannen rör basen samtidigt
En kvinna viker tvätt på golvet framför en rekyl.
En surfare som hoppar en våg på en surfbräda.
En surfare får luft medan andra tittar.
En manlig cyklist drar före flocken med grå, vit och röd ridutrustning, hjälm och solglasögon.
Hästen hoppar över hindret när en publik tittar på.
Två unga män möter varandra med medeltida rustningar, vapen och kläder.
En person hugger lök i en skärare.
En kvinna i bikini nedredelen håller upp sin högra hand nära en boll.
En man i grå t-shirt jonglerar bowlingpinnar.
En ung kvinna sitter på en grupp stolar medan hon poserar en blick.
Den unga damen skar gärna färska grönsaker till sin middag.
Sex personer i mid-evil stil kostymer bär styltor av varierande längd passerar av en grupp åskådare.
Två män i militäruniform står vid ett räcke medan en talar i telefon.
En mycket man på en motorcykel och två män på en vagn reser ner för en dammig två körfältsväg.
En man spelar ett tv-spel.
Flera cyklister på en stenväg, med åskådare tittar.
Folk gör köer för att göra sitt köp i antikaffären.
Två vita hipsters hanar slår varandra med kuddar på en offentlig utomhus torg.
En baseballspelare har gjort en intensiv pjäs för att komma till en bas, medan försvararen har förlorat sin balans.
En liten pojke som gråter bredvid en myntdriven åktur.
Två personer kör motorcykel i ett lopp.
En kille som heter Peter sätter upp något bakom en miniatyrjärnväg och andra människor i ryggen tittar på något på en drop-down skärm.
En massa motorcykel racers i färgglada hjälmar racing hals till hals.
En kvinna med brunt hår målar en bild på en staffl medan hon sitter ute.
En man håller i en stor vattenslang medan en annan man tittar.
Två män och en kvinna inspekterar framdäcket på en cykel.
Fem personer tävlar mot varandra med gokart.
Två personer som kör blå och svarta go-carts kör bredvid varandra.
En kock från Hodo Soy häller smet i en skål.
Två kvinnor, den ena håller i en sked och den andra håller i en plastflaska, lagar mat vid ett tillfälle.
En dam och en gentleman som bär blå handskar lägger något i en blå mugg.
En man som bär en trådlös mikrofon ler när han står nära en TV - skärm.
Tre flickor som andas in rök av något slag.
En man i blå uniform som sparkar en gul fotbollsboll med en nikeskylt på.
En bred uppvisning i finalen.
En fjäril har landat på huvudet på en blond liten pojke.
En pensionär i en sjukhussäng.
En grupp män som spelar fotboll, de flesta tittar på en man i svart.
Lilla flicka i gul skjorta sippar en bitter smakdryck.
En ung asiatisk man och kvinna står öppen mun framför mikrofoner, de är klädda i rockabilly stil och mannen har en blå gitarr
En svart hund står på en klippa, gröna fält bakom honom.
Ett litet barn som bär hatt leker på stenar vid kanten av en vattenförekomst.
En rugbyspelare i en vit och röd jersey skakar en tackling från en medlem i det motsatta blå laget.
Rugby spelare spelar ett intensivt spel av rugby, där bäraren hanteras av en medlem av det motsatta laget.
En man kajaker i en blå och vit kajak genom forsar.
En äldre kvinna smeker ingefära ett barn och håller honom mjukt för att lugna barnet.
En man med topphatt har en stor mugg på en pub.
Två kvinnor tittar på en kamera, en är kortare med brunt hår, medan den andra är blond och lite längre.
En liten pojke i en pool.
En kvinna i ett rött förkläde ger sig i väg mot ett urval av olika brödkakor bakom sig.
En man hukar sig ner för att ta en bild.
Pojken ser bakåt på kameran medan han rider i en gunga på en nöjespark.
En person i ett rum tänder en cigarett medan han håller i en katt.
En skallig militär i kamouflagekläder och ljusblå handskar knäcker ett ägg i en skål av rostfritt stål.
Tjej i röd outfit hoppar ur däck sving
Två män framför ett stycke musik, den ena i en rutig skjorta som sjunger in i en mikrofon och den andra i allt svart smetande en akustisk gitarr.
En lockig liten flicka ligger på stranden och tittar ner på vattnet.
En blondhårig pojke, klädd i blåmönstrade shorts, springer genom vattnet, som en våg avtar.
En fotograf tar en bild av ett lag som bär rött.
En ung hane går för en lek med en annan försvarar honom i en match av en-mot-en basketboll.
Barnen jagar en stor bubbla runt gångvägen.
Ett fotbollslag står på planen och väntar på sin tid att göra ett drag.
Tre fotbollsspelare kämpar för att få bollen.
En person på en parasail hoppar av en våg.
Två unga fotbollsspelare tävlar om bollen.
En grupp på 5 unga flickor poserar för ett fotografi genom att försöka hoppa i luften precis som bilden tas, en av dem stannar på marken och håller en spädbarnshane.
Två barn springer längs en trottoar klädd i kostymer.
Två personer tävlar i ett rullstolslopp på en stadsgata.
En man i kostym har vatten.
En man som försöker binda en liten ko med ett rep.
En kvinna i röd skjorta och lila hatt bär en blå behållare full av föremål på huvudet.
En man som bär en blå hattsten klättrar upp för ett brant rockansikte.
Tillsammans med medlemmar i det lokala hockeylaget går en beslutsam kvinna den sista sträckan mot mållinjen för maraton.
En kvinnlig löpare klädd i en sporttank och kort hejas på av en skara åskådare.
Ett par förbereder för avfärd i sin yacht.
En domare i en roller derby tittar på kvinnliga åkare när de passerar förbi.
En man som kastas i luften medan han trampas ner av en tjur.
Två soldater tränar en polishund när den hotfullt tar tag i ett av soldatens träningsredskap med munnen.
Mörk bild av män spela bongo trummor och dricka
En första baseman i en dams softball spel försöker tagga ut löparen i slutet av en pickoff spel.
En man som vindsurfar i havet.
Fyra barn leker vid en fontän utomhus.
En kvinna målar en scen av Grand Canyon på sin bärbara staffl.
En barfota man fotograferar ett par som ligger i det gröna gräset under några palmer med vatten.
En grupp äldre tittar på en föreställning.
Fyra tjejer spelar fotboll på ett plan när deras tränare tittar på.
En söt ung pojke som viftar med en amerikansk flagga utanför.
En tonåring utför ett trick hoppa på en stad gatan hörnet.
En ung kvinna i lila löparskjortor rider en röd cykel i staden.
En hona i en gul badmössa simmar i en pool.
En skjortlös man framför en uttorkad tegelvägg utanför.
En ung flicka i en skara människor som snurrar två hulahoops på en gång.
En ung vit man i löputrustning joggar vid vattnet.
En man med ett ben som kastar diskusen.
Denna version av street hockey är på mellan organiserade lag.
Människan höjer sina armar triumferande som han leder flocken i en cykel tävling.
Små barn har en rolig sommardag genom att leka i vatten.
En manlig skateboardåkare åker av stegen för att göra ett trick drag för kameran.
Pojken slickar glasyren från skeden.
Männen är mycket påhittiga och lyckades till och med ta en tupplur även i detta ovänliga utrymme.
En fotbollsspelare i luften när han sparkar fotbollen.
Någon rycker nerför en hög klippa med solen och molnen på himlen.
Manlig publik surfar på en konsert.
En domstol-sidan action skott av flera professionella basketspelare i ett spel.
Två män spelar gitarr medan en kvinna tittar bakom dem.
En man som bär en blå skjorta talar i mikrofoner mitt i en bakgrund av tecken.
Två unga kvinnor i färgglada kläder går genom våtmark.
En flock hästar stänger ihop precis utanför grinden vid en hästkapplöpning.
Två män som tittar på varandra och spelar pool.
En grupp hästar och deras jockeys tävlar över gräset.
Surfaren hukar sig lågt och rider vågen.
En man gör en vända medan en publik tittar.
En fotbollsspelare springer förbi sin tävling med bollen.
Fem män som står på en musikscen ler och vinkar åt en osynlig publik.
En kille i vit t-shirt på en Mac-dator.
En lång äldste man står med sin hand runt en annan kortare äldsteman mitt i staden
En DJ värd tar micken och samlar sin publik.
Ett gäng löpare hoppar över ett hinder, och två av dem faller i vattnet under det.
Brunettkillen är klar med ett hopp i valvet.
En hög hoppare är mitt i hoppet medan hon fortfarande håller i stången.
Två fotbollsspelare är på planen framför en stor publik.
En man springer, i en gul löpare skjorta och matchande löparshorts, längs vattnet med en stor stad i bakgrunden en vacker dag.
En motorcykelåkare färdas längs en lång grusväg kantad av gröna träd.
En stor fotbollsspelare tar itu med och tar ner en annan spelare från det motsatta laget mitt i ett actionpackat spel.
En muskulös muskulös man petar bröstet med en brun dolk medan han grimakerar.
Ett lag av fotbollsspelare alla klädda i vitt och grönt två av dessa manliga spelare tittar på en telefon leende.
En man i en unik kostym spelar säckpipa medan vissa stirrar på honom.
En långhårig man i en blå skjorta jonglerar med sex apelsinbollar.
En man, med glasögon och en vit skjorta, radar upp en biljardbild.
En grupp människor står i kö längs ett svart staket.
Mannen tittar på motorn i den gamla brandbilen.
En man i blått intervjuar en man i mörk kostym medan han sitter i ett vitt tält.
En vuxen och två barn leker i högar av fallna löv.
En kvinna och en man skar ihop degen i små bitar.
En liten pojke som leker i sanden på stranden.
Två barn leker med sand på en strand nära havet.
En grupp människor gräver hål i jorden.
Två krigsartister slåss inför en grupp människor.
Tre soldater försöker släcka en brand med en brandslang.
En kvinna med lila skjorta och vit hjälm rider en brun häst.
En vackert klädd liten flicka poserar i skogen med sin promenad käpp.
En kvinna håller en drink i ena handen och pekar på en målning med den andra.
Tre killar som spelar golf längs en vattensamling.
En kvinna går längs stranden med tre barn som följer efter henne.
Detta visar många människor på cyklar i olika färger uniformer och hjälmar.
En man sitter vid en datorstation bredvid en kvinna och använder datorn.
En medelålders solomusiker uppträder genom att sjunga och spela gitarr.
Med en fasad i bakgrunden står en man på en annans axlar och håller flera brinnande pinnar.
En ung pojke som gör sig redo för en fiskedag.
En man i svart baddräkt spelar volleyboll på en strand med palmer.
En kille som sitter i en stol rakar sig.
Några personer på en båt med ett vitt hus i bakgrunden.
En cyklist racing i ett cykellopp.
Grupp av personer som står framför en affär som säljer cyklar för barn.
En pojke, med blå glasögon, simmar i en pool.
En kvinna övar sin form med ryggsim under varv simning vid en lokal inomhuspool.
Två män och en kvinna spelar musik på en scen.
Två kvinnor i lila glänsande klänningar dansar framför buskar.
Fyra vuxna som spelar baseball, med en skog i bakgrunden.
Kvinna tennisspelare i en grön och röd klänning balanserar en boll på racket.
En man som försöker nå tennisbollen i ett tennisspel.
Flera killar spelar cricket på ett plan, medan en gammal man och dam tittar i bakgrunden.
En grupp människor på en brygga vid en stad som går ombord på olika båtar
En bebis med brunt hår i flätor som sluter ögonen.
En smedja förberedde sina verktyg i sin enkla verkstad.
En grupp pojkar tittar på en pojke klädd i svart med blå strumpor sparkar en fotboll i luften på sanden.
Två dansare i rosa toppar och randiga capri bottnar uppträder på scen barfota.
Två vita hundar leker på gräset.
Hmong mamma tvättar sina barns kläder med vacker natur bakom sig.
Närbild av en militär man och kvinna i en blå klänning som dansar på en militärbal.
Fyra barn ritar bilder på en stor vit duk.
Människor står och sitter vid runda bord i ett stort rum.
Fem små flickor poserar i matchande danskläder.
En målning av människor som står utanför byggnaden under två träd och ser mot ett gult ljus.
Man med röd rock och spetsigt hår blåser på en kazoo på scenen.
En ung man surfar på vågens krön.
En person är kitesurfing vid en bro.
En man som håller i en kamera sträcker sig över ett räcke för att skaka hand med en examen från 2012.
En medelålders man och kvinnor i en blå skjorta tittar på mannens diplom.
Förutom en tegelbyggnad kramar en kvinna en nyutexaminerad i gratulationer.
I ett urbant område agerar människor ut sitt dagliga liv genom att gå, äta och njuta av sällskap.
En man träffade precis bollen på golfbanan.
En grupp artister klappar på scenen.
Folk i bakgrunden sitter och ser på när två flickor i röda skjortor gör volter.
En grupp hejaklacksledare utför stunts på ett spår.
En ung kvinna i en prickig skjorta och glasögon framför några träd.
Två barn fotbollsspelare brottas för bollen.
En äventyrlig skidåkare rörde sig skickligt nerför den branta, snöiga sluttningen med hög hastighet.
Runners jogging genom vatten med en regnbåge visas.
Den ene är skjortlös medan de andra två arbetar med att bygga.
En asiatisk man i militären gör armhävningar för en överordnad.
En ung flicka med rosa tärningar i sitt bruna hår har en sorglig blick i ansiktet.
En man försöker fixa ett färgglatt föremål.
Den lille pojken går nerför trottoaren i sina mammors skor.
Två personer som leker med en volleyboll i en pool.
Två fotbollsspelare, en klädd i vitt och en klädd i blått, rycker varandra samtidigt sparkar rosa och vita bollar.
En fotbollsspelare jagar en boll mot en sidolinje på planen.
Två fotbollsspelare jagar en medlem av motståndarlaget som försöker få kontroll över bollen
När konfetti flyger, firar ett fotbollslag i vita uniformer.
En våt brun hund hoppar upp för att få en vit basketboll.
En tjej med auburn-hår sitter vid ett bord och tittar över axeln.
En man tävlar om ett cykellopp medan de andra cyklisterna är direkt bakom honom.
Män, kvinnor och barn samlas runt med spadar plocka upp stenar.
Mannen, utan skjorta, sträcker sig i en hink för att utvinna ämnet inuti.
En ung mor och hennes barn går längs en gata.
En grupp ungdomar som samtalar lyssnar på när de håller i en drink.
Två vita kvinnor som har ett samtal och en öppen öl.
En man som håller i en påse ger en annan man en grisryggfärd framför en sandwichbutik.
En man och en kvinna dansar lyckligt.
En flicka som håller en uppstoppad Psyduck leksak ler medan hon sitter på en säng.
Barn leker i fontäner som sprutar vatten från marken.
Män i ett cykellopp går nerför en kulle
Ett band, bestående av minst en manlig gitarrist och en kvinnlig sångare, spelar musik på en scen.
En kanna och catcher på ett baseballfält med bollen i mellan dem.
Violinsolister tar scenen under orkesterns öppningsshow på teatern.
En man som springer i ett maratonlopp springer över en bro.
Två livräddare vakar över havet en molnig dag och en amerikansk flagga hänger bakom dem.
En man som sitter på trappan med ett barn som åskådare går förbi.
Ett leende barn som ger sina föräldrar en färgglad godbit.
Fyra bicyklister som bär hjälm tävlar längs en stadsgata medan åskådarna observerar.
En cyklist rider en gul cykel med ett fält i bakgrunden.
En ung pojke och flicka dras i en barnvagn dekorerad som den amerikanska flaggan.
En ung pojke leker med sin boll framför en byggnad.
En ung flicka, som bär en gul tanktopp, leker utomhus med andra barn i bakgrunden.
En konstnär ritar en karikatyr från ett fotografi, bredvid honom finns flera kändisteckningar.
En grupp män kör en street race medans de bär idrottsutrustning och sina racer nummer.
Marathonlöpare som springer mot mållinjen.
På en liten flod drar fyra rödklädda roddare sin gula båt framför flera andra.
En brottningsmatch pågår medan en publik tittar.
Två män som övervakas av många, utan byxor eller skjorta, en som har tatueringar och bär någon form av huvudbonader.
Två män i separata kajaker genom forsar.
En pojke som hänger upp och ner på en stege bredvid en annan pojke som klättrar upp i ett knutet rep.
Två män boxas utan tröja med svarta byxor på
Två blonda barn, en pojke och en flicka, håller käppar och ler.
Två vänner tävlar i ett tävlingslopp.
En man skjuter en pistol utomhus, på vad som ser ut som en vacker solig dag.
En kvinna med brunt hår och marinblå jersey springer
En kvinna springer på ett tävlingslopp och håller i en flaska vatten.
Tre vita män sjunger och uppträder på scen på en konsert.
En svetsare som bär en svetsdräkt är svetsskrot tillsammans.
Att spela teeboll är så kul för den här lilla pojken.
Två kvinnor tävlar i ett maraton, medan en liten pojke tävlar nära bakom dem.
Män och kvinnor på scenen håller stolpar med färger och utför.
En tjej i en röd tank topp pratar på en mobiltelefon.
En kille som ligger på ett fält som verkar väldigt lycklig
En man håller ett litet barn på en trädlem.
Fem musiker som håller sina instrument poserar för ett foto framför en bakgrundsbelyst båge.
Fem musiker, tre kvinnor och två män som ser ut över en vägg med sina instrument bakom ryggen.
Fem personer bär svarta och håller musikinstrument tittar uppåt.
En kvinna i rutig klänning och bara fötter utför en rituell dans över bambupålar.
Ryggen på en persons huvud visas, när de kliar huvudet med handen.
En man klädd i orange och svart kör ett maraton genom gatorna när folk tittar på.
En grupp löpare tävlar i ett sommarevenemang.
En simmares hand tas när han kommer upp ur vattnet.
Flera män i våtdräkter och glasögon som står bakom ett band.
En stor grupp simmare i våtdräkter och badmössor dyker ivrigt ner i vattnet.
Ung kvinna njuter av att spela pool.
En liten flicka på ett baseballfält som svänger på en baseball på en tee.
En ung kvinna hoppar i luften på en skateboard.
Ett barn med dreadlocks breakdansar på en offentlig trottoar.
Sanitetsarbetare på lovet mitt på dagen.
En man använder en slägga för att hamra en ring på en tunna.
En kvinna som bär en röd jacka på gatan.
En brun häst med vit man gör ett trick med en man som sitter på ett fält.
Tre personer från ett land i öster dansar på ett dansgolv.
Tre män i militärdräkt som gräver sand i en öken.
En uniformerad officer talar in i en kommunikationsapparat medan han sitter.
En man som bär armékamouflage står bakom ratten på det fordon han opererar.
Person som flyger i luft med sandaler, glasögon och vinddräkt.
En gitarrist uppträder under en konsert tillsammans med sin bandkamrat, på basgitarr.
Tre unga vuxna diskar i köket.
En kvinna i svarta shorts och en lila topp, jogging medan du trycker på en grå barnvagn med ett litet barn i barnvagnen.
Kvinnan i blå huvudduk och svarta kläder bär 2 brickor bakverk utanför en byggnad.
Tre unga mörkhyade män sitter på staplad frukt och ler mot kameran.
Utomfältaren dyker för att fånga popupen på mittfältet.
En fotbollsspelare följer igenom med en spark som en andra spelare klockor.
En person breakdancing medan några unga pojkar tittar.
Folk tittar på en ung pojke som ser ut som om han faller ner på botten på ett kaklat golv.
En man i glas som arbetar med en matberedare och står bakom ägg, mjöl, apelsiner och smör.
En brandman klättrar upp för en brandbilsstege.
Två män med blå fotboll uniformer tränar fotboll.
Barn som bär hattar och gör roliga ansikten medan de ler står bredvid ett staket i sanden.
Killen i röd uniform studsar en fotboll av huvudet.
Två fotbollsspelare springer och sparkar en fotboll på en match.
En kvinna är i vattnet redo för wakeboard.
Två kvinnor som spelar badminton med träd i bakgrunden.
En flicka med orange väst rider en brun häst.
En ung man i svart hatt och vit t-shirt är upphängd i luften på sin skateboard.
En racerbil driver på den obelastade vägen.
En aktiebil tävlar längs en grusväg och sprutar en plym av smuts bakom den.
En förare kör för fort en liten bil mycket snabbt.
En pojke i svart hjälm hoppar en cykel med en liten stad synlig i bakgrunden.
En kvinna med glasögon och en läpp piercing sitter ner tittar på sin rosa iPhone.
En man spelar på en stand up bas genom att plocka strängarna.
En mamma tränar i en vacker trädgård.
En person bär en liten kajak eller båt till vattnet medan två andra tittar.
En flicka skriver på sin dagbok på en picknickduk.
Tre stadsarbetare i hårda hattar häller cement från en lastbil och lägger trottoaren.
En baseballspelare som är på väg att ta en inkommande baseball.
En man som visar sin akrobatiska skicklighet med en monoboard bogseras bakom en båt på en sjö.
En sångare i vit rock som sjunger in i mikrofonen.
Ett tecken med ordet försäkring skrivet i rött är fäst vid en stolpe.
En äldre svart man som använder en symaskin på en skjorta.
En kvinna i rock drar sin utvalda tall genom snön.
Pitcher på pitching hög i maroon keps och jersey släpper baseball.
Två pojkar vilar på en stock som flyter längs stranden av en vattensamling.
En baseballspelare vid University of South Carolina som slog en boll med ett slagträ.
En man i svarta kläder rider en ATV längs en väg.
En person med vit och svart kostymbräda som vaknar upp i vågorna.
Två unga flickor som bär vita tennisuniformer skakar hand.
En broder som håller sin yngre bror ute i kall luft.
Ung pojke i en blå och grå tröja som håller en trästolpe.
Vissa män lär sig kampsport.
En grupp män ser två män uppträda på ett gräsfält i ett område.
En grupp vuxna och barn med en vit elefantstaty på en festival.
Fyra män i mångfärgade löparkläder och skor sprintar nerför en gata medan åskådare titta.
En man i vitt organiserar en gul mapp.
En pojke i svart och grön t-shirt som leker utomhus i sanden.
En man med glasögon håller ett mycket ungt spädbarn.
En tubaspelare klädd i formell klädsel uppträder tillsammans med sina bandkamrater, en banjospelare och en trumpetspelare.
En kvinna med en svart skjorta på grillar kabober.
En kvinna tvättar en skål framför ett fönster med nyanserna dragna.
En rödärmad man har kastat ner, på ett sparrande sätt, en gentleman med blå ärmar.
En byggnadsarbetare står på en kran och lägger en stor arm ovanpå en ställning som pågår.
Ett fotbollslag springer när sparkaren rör fotbollen med foten.
Två män tävlar om bollen i en fotbollsmatch.
En fotbollsmålvakt hoppar upp för att rädda bollen från att gå i nätet.
En man i fotbollsuniform sparkar bollen medan en annan man tittar i bakgrunden.
En person flyger genom luften i ett fält på en motoriserad smutscykel.
En dam i glittrig klänning spelar gitarr och sjunger in i en mikrofon.
En grupp barn som går på en stig.
En man i röd skjorta som rider på en häst i vad som verkar vara en rodeo.
Två oentusiastiska barn sitter i en parkerad brandbil.
En stadsarbetare (med orange väst) som arbetar på en bärbar dator som sitter ute på marken.
En kvinna som bär solglasögon rider en brun häst.
En motorcyklist flyger genom luften ovanför en grusväg.
En man i vit skjorta och rutiga shorts sätter sig ner.
Målvakten vänder sig om för att se pucken i nätet, medan laget stiger från bänken.
Två hockeyspelare åker skridskor på isen.
Person som bär cowboykläder kastas av en tjur medan han omges av rodeo åskådare.
Man på häst bär vit hatt försöker lasso lilla djur.
En naken bebis och ett litet barn smetar varandra i färg.
3 män, 2 skyfflar smuts och den andra lägger ner cement.
En man som surfar på en våg med några personer bakom sig som simmar.
En surfare som rider på en våg i det blå vattnet.
En manlig surfbräda i svart våtdräkt rider en enorm våg i vackert blått vatten.
Två kvinnor sitter och spelar på ett kasino.
Två barn sitter utan tröja på en studsmatta.
En asiatisk kvinna har en liten flicka.
En man i randig skjorta hoppar från en gunga.
En man lagar en ostburgare till en kund.
En man sparkar en annan man i huvudet i en röd ring medan en annan man tittar.
En flicka som står utanför en klädaffär
Två bulldozers transporteras på en lastbil med träd i bakgrunden.
Kvinna försöker slutföra en reserv i bowling med hjälp av en röd boll.
En kvinnlig dansare poserar på tå i en elegant fotostudio.
En man fäster cyklar på baksidan av sin bil på en trädfodrad parkeringsplats.
En brun och vit hund som springer med tungan hängande ut.
Två människor går sina hundar på stranden, med en molnig himmel.
En skoputsande man sitter på sin pall framför en tom stol.
Två män slåss med en spade och toppen av en grill.
En person i en ljusblå outfit tävlar en smutscykel genom en kurs i skogen.
En grupp skolbarn som tittar på en grupp män som bär vita skjortor
Två män skakar hand utomhus framför flaggorna
Mamma försöker ändra roll med sin son i köket.
Turister, båda kvinnor (en äldre, den andra betydligt yngre) poserar med låtsasastronaut för bild.
En man leder en orkester när alla andra musiker följer hans ledning.
Människor som omger ett teleskop för att se saker och ting på långt avstånd.
En kvinna som sjunger i en klubb med glasögon och spelar tangentbord
Två gamla män sitter i en bubbelpool.
Två flickor går längs en stock på ett fält utanför.
En man med ett stort nät står i vatten som är upp till bröstet.
Hästar och jockeyer springer i en turf race.
En Jockey i blå hjälm, röd skjorta och vita byxor rider en tävlingshäst med "sparkasse" skyltar i bakgrunden.
Två män brottas mitt i höga byggnader.
En gitarrist, en trumpetspelare och två saxofonister tar scenen.
Två män i havet surfar på brädorna och försöker fånga vågor.
Tre personer paddlar kajak och två har kraschat in i varandra.
Två kvinnor utsmyckade i traditionella stamkläder står utanför.
Man klädd i svart kör dramatiskt en racing motorcykel längs en sträcka av gatan trottoaren.
Två racerförare i en liten racerbil med åskådare i bakgrunden.
En skäggig man med blå skjorta och vit t-shirt arbetar på ett fiskenät.
En liten pojke i orange kragetröja svingar ett basebollträ.
En vandrare klättrar över klippor för att komma närmare ett vattenfall i ett landsbygdsområde.
Cowboys kämpar för att krångla hästar på en arena som åskådare tittar på från läktarna.
Cykelhjul i förgrunden med några män i jackor suddigt i avståndet.
Två asiatiska kvinnor dansar och bär färggranna kläder.
Ett litet barn, som bär hjälm, rider en BMX cykel på en grusväg.
Två män inspekterar den yngre pojkens arm för skador.
En grupp människor samlas och i mitten tar en kvinna sin hand till en mans ansikte.
Män och kvinnor dansar tillsammans i formella kläder.
Ett gäng barn i gula hattar tittar över ett stängsel.
En dam och en ung pojke är under paraplyet.
En motorcykel racer tar en kurva på en gata krets.
Tre personer skyfflar sand.
En man i gul och svart våtdräkt surfar på en liten våg.
En svart man som tittar och sträcker armarna uppåt.
Tre män med öronskydd håller i en pistol och övar på att skjuta på skjutavstånd.
En man med blont hår och glasögon spelar en typ av horn.
En äldre herre bär en tikilampa nerför en gata kantad av människor, eftersom några av dem fotograferar.
En man illustrerar med hjälp av en sprayburk.
En svart man spelar gitarr medan en kvinna i en mörkgrön rock i närheten tittar bort.
En rodeospelare tas ner av en tjur.
En liten pojke som leker i klippor och sand nere vid vattnet.
En grupp infödingar samlas i en infödingsbutik.
En baseballspelare i vitt förbereder sig för att kasta bollen.
En baseballspelare slår bollen som en huk bakom sig.
Två barn har grävt ett stort hål vid stranden och fyller det med vatten.
En pojke skyfflar sand på en strand.
En flicka, som knäböjer på sanden med en rosa Minny Pigg hink nära henne, kastar en skopa sand med en spade.
En man i röd kostym utför motorcykel stunts.
Ett dussin fotbollsspelare i svarta uniformer står i en rad på ett gräsfält, deras andetag synliga i den kalla luften.
Tre unga killar som jobbar i ett mörkt rum.
Man i en blå motocross outfit och röd hjälm rider en smuts cykel på ett spår.
En äldre man håller en hammare medan han tittar på något vi inte kan se.
En gitarrist, en trummis och en annan bandmedlem uppträder på scenen med rött ljus på bakgrunden.
Barn njuter av en åktur på en karneval.
Tre män i ett rockband som uppträder på scen, i hög modekläder och långt hår.
Männens roddlag i deras gröna båt övar för sin kommande säsong.
Två personer på cykel racing på banan rundar ett hörn
Två män på motorcyklar tar en sväng på ett spår.
En blek vit dam med blont hår och kristallklara blå ögon, somerly poserar med två röda bär placerade i hennes näsborrar.
Man surfar ombord med sin hund i havet.
Sju män med byggnadshjälmar arbetar på järnvägsspåret.
Två personer ro en båt när en flock fåglar passerar dem.
En grupp båtfolk som seglar på en slingrande vattenväg.
En man åker skidor i vatten.
En svarthårig man sover på en bänk på en gata.
En man med en handtruck tittar på gul graffiti.
Köksmästare lagar mat utomhus med bröd och matlagningsutrustning synlig bredvid de ingredienser de arbetar med.
Tre åskådare ser en joggare passera när en av dem ger honom en drink.
Två män, en i en röd jersey med en boll och den andra i en blå jersey, springer på ett gräsigt fält.
Män klädda i militärkläder övar sina rundor.
En skiplastare flyttar smuts i en skog medan 2 män tittar och direkt.
En man som går på smuts på en byggarbetsplats.
Två män arbetar hårt i det som verkar vara snöröjning.
En dam skriver på en tavla.
Två äldre kvinnor spinner trådar på snurrande hjul, klädda i gamla kläder.
En kvinna i vit klänning som håller blommor stående framför 4 kor.
En pojke med röd hatt står mitt på vägen.
Två män står på däck på ett stort skepp
Två män, klädda i hårda hattar och blå och gula rockar står framför en stor maskin och ler.
Två män står i en öppen dörr till en galge, med den tredje mannen inuti.
Ett asiatiskt barn som är klädd i rött gråter som en asiatisk kvinna verkar trösta henne.
Två lag spelar fotboll i en stor stadion som är fylld med åskådare.
En ung dam utför yoga tillsammans med resten av sin klass.
En man klädd i kamouflagefärg håller i en pistol och riktar den mot sitt mål.
Två män i vitt övar fäktning på en domstol.
En skateboardåkare landar ett trick från en hög plats.
En bartender i svart skjorta förbereder en rosa drink i ett martiniglas.
Tre personer på cyklar i startlinjen av ett lopp.
En liten pojke och en liten flicka bär formella kläder på ett bröllop, medan de går nerför gången.
En cykelmekaniker förklarar fysiken hos en cykel till en registrerad sjuksköterska.
En indisk kvinna som sitter ner med handen utsträckt, i en blå klänning och dyra smycken.
Låt oss se hur många människor vi kan få att stirra på oss.
En man på scenen som pratar genom en mikrofon i en svart skinnjacka.
Javelin kastare bär en mörk skjorta och förbereder sig för att kasta.
En vitklädd ryttare på toppen en häst hoppar över en rad stolpar.
En person rider en vit häst medan han hoppar hinder.
En kvinna med blå stövlar som står framför en stor korg med grönsaker.
En lockig man i kostym spelar trumpet i sidled.
Arkeologer gräver efter nåt.
En enda person som cyklar.
Två personer rider cyklar bredvid varandra på marken med gräs i bakgrunden.
En kvinna i vit skjorta och shorts spelar en röd gitarr.
En liten pojke håller en tänd glittrande i trädgården.
En racing katamaran skär genom vattnet.
En katamaran på havet i en seglingstävling.
En grupp vänner gör sig redo att gå på ett vattenäventyr.
En tjej i en grön tröja topp och blå shorts gör sig redo att sparka fotboll nära målet.
En gammal flintskallig vit man äter en liten tjejkex.
En man som kör på gatorna med en cello i en huvtröja och ryggsäck.
En kvinnlig softballspelare som svänger på en softball.
En ung flicka som bär en röd skjorta med höger arm upphöjd och vänster arm har en softball handske.
En liten pojke sitter i en gunga.
En skäggig man spelar flöjt, och en person med fasor som står bakom honom spelar ett annat instrument.
En man i vit skjorta och keps bakar kakor.
Ett barn med gröna hörlurar på vinkar åt en stor skara människor.
En arméhund som tränas av en soldat.
En kvinna i svart förkläde står framför en spegel.
En man som bär glasögon simmar i en pool.
En vit hund kommer fram från en gul tub på en hinderbana.
Den unga flickan är rullskridskor utanför nära gröna buskar.
Tjejen i det vita basketlaget high-fives en medlem i det svarta laget, medan andra tjejer samlas.
En flicka står på en pire när en färja kommer in.
Kvinnor i svart klänning tar bilder av barn framför blommor.
Ung skateboardkille vänder på sin bräda medan han utför ett stunt.
En man bär många väskor fyllda med föremål när han ler mot kameran.
Fyra personer på en semesterfest på natten.
En man cyklar på en liten bro över en vattensamling, kanske ett träsk.
En italiensk idrottsman poserar på planen.
En liten utställningshund sprang bara genom ett orange flexibelt rör.
En leende kvinna med slutna ögon svingar på en däcksvinge.
En ung pojke i gul skjorta drar med en blå krita vid ett litet utfällt bord.
En liten pojke med blont hår sitter på golvet och klipper något med sax.
Två män spelar backgammon medan en tredje tittar på en trottoar.
En ung pojke är i ett överväxt fält med en leksak gräsklippare.
En scen med en stor skärm och en publik på cirka 100 personer.
Det finns en tätbefolkad strand med klart vatten.
Hunden sticker ut tungan och går i gräset.
Tre segelbåtar i ett seglingslopp.
En kvinna i randig skjorta använder en skärbräda och knivar för att skära några grönsaker.
En man och en kvinna som står framför en svart stationsvagn.
En kvinna i en kort, ärmlös ljus orange klänning och svarta leggings sitter på en cement bänk tittar ner, med många cyklar parkerade bakom henne.
En cyklist i röd uniform avrundar en kurva på sin cykel.
En äldre man bär den olympiska facklan för OS i London 2012 förbi en grupp åskådare.
En man i olympiska kläder bär London 2012 facklan ner på en gata.
Tre människor ler när de väntar på att deras ras ska börja.
En pöbelhop har samlats i protest; en kvinna bär ett tecken på hebreiska.
En akrobathona som bär en röd och vit randig skjorta och blå byxor uppträder på en stolpe.
Man håller en kopp och toalettborste bredvid en urinoar.
En man i blå skjorta pratar på en mikrofon, framför folk som sitter ner.
En man i hjälm som cyklar.
Två män målar graffiti på en vägg.
Asiatisk man i rött och svart spelar basket.
En man med svarta byxor och hjälm rider en brun häst.
Föräldrar engagerar sig i utomhusmusikfestligheterna genom att hjälpa barnen att spela handfat.
En kvinna står bredvid en målning hon kan ha målat.
En hona sjunger in i en mikrofon under en utomhusrockbandskonsert.
En professor framför sin klass håller en föreläsning.
Det finns fyra män, tre sittande och en stående, bär samma mörkblå uniform.
En clown leker i en park med bubblor, medan ett litet barn leker.
En cyklist i rött knuffar sin cykel.
En gammal, kanske hemlös, man sitter vid ett bord med ett glas framför sig.
Folk i kostymer väntar på att uppträda på ett evenemang.
En man i vit skjorta sitter på mobilen vid grinden.
Motorcykelpolis rider i en parad.
Två män i röda skjortor står med en man i svart skjorta.
En man maler sin skateboard på ett skyddsräcke.
En kvinna deltar i en träningskurs med kickboxing-stil rörelser.
En ung pojke med grön väska står bakom en stolpe i en tunnelbanestation.
En kvinna spelar bas och sjunger med sin bandkamrat med är en man som spelar gitarr och trummisen spelar i bakgrunden.
Den lilla pojken springer och ler.
En man klädd i vitt med guldränder som håller i en gyllene fackla som viftar mot folkmassan.
En äldre man på ett politiskt möte med en skylt som tackar våra trupper.
Personen som kör en "en man" sätter den på två hjul i sanden.
En man rider en ATV genom öknen.
En dune buggy med en manlig passagerare får lite luft när den kör över en sanddyn.
En erfaren fyrhjuling som skyndar på några sanddyner.
En asiatisk man bär en kimono medan han övar sin kampsport med en kollega.
En ung skolflicka ler mot kameran.
En grupp barn på en karusell och lekte i parken.
En grupp människor som spelar karnevalspel.
Profil vy över en man med en brun pipa i munnen.
En liten pojke som ler och rider i en spade.
En liten flicka har doppat huvudet i en skål med vatten.
Kannan kastar bollen i en basebollmatch.
Den #5 basebollspelare från Green Team försöker göra fånga som #7 Gray Team spelare korsar basen, med umpire tittar på att göra samtalet.
En man leker med ett barn och håller upp honom i luften.
Två tjejer och en kille är inblandade i en pajätande tävling.
En korthårig man hoppar på ett stort stenblock.
I vad som verkar vara en patriotisk parad, en man som rider ett fordon håller en liten flicka och amerikanska flaggor i överflöd.
Män som bär förkläden, hattar och solglasögon grillar.
En grupp människor sitter vid ett långt bord med vinglas.
En ung pojke som stänker en äldre person med en flaska vatten
En man och en kvinna spelar alla akustiska gitarrer på scenen, omgivna av högtalare och mikrofoner.
En vuxen man i kamouflage hjälper ett litet barn att hålla ett gevär.
En man som syr ett plagg med en antik symaskin.
Ett barn sprutas med vatten medan äldre människor sitter och tittar.
En man och en kvinna åker skridskor på en rink.
Tre män i hårda hattar styr stora maskiner.
Ett ungt par sitter i en roll och äter glass när barnen leker och andra har kul omkring sig.
Folk njuter av avkoppling och läsning i denna gröna och skuggiga plats.
Ung man på en surfbräda rider en tuff våg.
Baseballspelare #38, Morse ses stående och tittar på kannan.
En man i gul skjorta fyller några tunnor med en liten scoop.
Två tjejer tittar ut genom fönstret på "Hair at Hart".
Bruce Springsteen, klädd i svart, håller i en mikrofon och pekar mot en publik.
En sittande man avfyrar ett vapen.
En bowlare har precis släppt en bowlingboll nerför gränden mot stiften.
En surfare som rider på toppen av en våg i havet.
En surfare surfar en stor våg på en vit surfbräda, bär en svart och röd body.
En man som surfar på en våg och hänger tio.
Det finns fem hästryggsryttare som rider genom en dal på en stig i solljuset
En kvinna och ett barn är på en fullsatt flygplats.
En fet polis och en fet dam sitter tillsammans medan polisen bläddrar igenom pappersarbetet.
En kille kastar vatten ur en blekhet i en fontän.
Många uniformerade cyklister går nerför en gata förbi bilar parkerade på sidan av vägen.
En kvinna och en ung flicka som klättrar upp på en gräsbevuxen kulle.
En liten pojke i ett leksaksrum som bär Batman pyjamas bygger något med leksaker.
En man med långt skägg som spelar gitarr.
En kvinna i en röd tank topp och en Men's Health hatt sitter på marken och äter sin lunch.
En brun och svart Yorkie leker med en röd boll.
En man tillverkar keramik och tittar noga på det föremål han gör.
En paintballer, duckar under en röd barriär.
Några av de tio barnen har juicelådor, en har en volleyboll.
Två män i orange skyddsvästar målar en trottoarvit.
Ett barn ser en man forma ett keramikföremål på en krukmakares hjul.
En kvinna som spelade fiol i en konsert.
Två män i solglasögon tittar på något framför dem.
En kille som lutar armen mot en stol med slutna ögon.
En afrikansk amerikansk basspelare som bär en blå skjorta och backas upp av en trummis.
Cyklare i antal rider ner i en parad.
Ett team av människor som lägger händerna i mitten.
En ung flicka som gör en backflow i vattnet.
En kvinna i bikini är i vattnet och hoppar i luften när hon håller i en zebraballong.
En kvinna som firade efter att hon bowlat en ram i en bowlinghall.
En mattjänstperson ger en kund sin dubbelscoopglass i en kon.
En bicyklist rider förbi som en publik tittar bakom en banner.
Två män i vita uniformer och blå hjälmar leker på ett bollplan.
En pojke slappnar av i en hängmatta vid en flod.
Ett barn står på en fotpall i ett kök vid köksdisken.
En manlig golfare försöker träffa golfbollen ur en sandfälla.
Ett fotbollslag firar en seger när en spelare hoppar på en annans rygg.
Ett band bestående av en hona och tre hanar spelar under dagen.
Två barn som bär solglasögon sitter utanför ett plasttält.
Tennisspelare i vitt svänger hennes racket.
En ung man är utanför och håller i en trådrulle.
Två bicyklister i ett lopp med hjälmar med åskådare i bakgrunden.
Man rider på cykel med vit och grön cykeltröja och hjälm.
Grabben är i vattnet och håller fast vid ett rör.
En simmare, med en blå mössa och blå glasögon, simmar i lugnt vatten.
Folk står och tittar på nån sorts samling.
En ung pojke klättrar i berg, medan han är upphängd i en sele.
En man tittar på ankor som hänger genom ett fönster i en etnisk mataffär.
Barn är alltid ett nöje att vara med och le.
En kvinna och en liten flicka tittar in i en utställningslåda.
Den ljusbruna hunden med vita fläckar nibblar på flickornas hand.
Unga flicka bär en bukett med blommor.
En familj på tre baskar i solen i en park.
Man rakar en annan mans ansikte med rak rakkniv.
En skjortlös man gräver bort sand med en rosa scoop medan en liten flicka tittar.
Killen gör rullskridskor och älskar det
En ung man i en grå huva och en blomma på huvudet slår en pose efter en måltid.
En hona snurrar i en vit klänning.
En folkmassa lutar sig mot barriärer längs en väg, medan en polis på en motorcykel kör förbi.
Mannen i gul skjorta håller i en mikrofon.
En man som bär badbyxor hoppar ner från en stor sten i en vattenförekomst.
En pojke simmar bröstsim på ett simmöte.
En blondhårig tjej som bär en mössa som blåser bubblor i en trädgård.
En grupp solbrända människor i en monter med grönsaker.
En kvinna sitter på ett konstverk.
En liten flicka i en röd regnhatt leker i leran med flera vuxna.
En grupp människor som städar några släktingar till havsdjur.
Män spelar basket inför en stor publik.
Två balettdansare, en klädd i vitt och en klädd i grönt, dansar på en scen.
En man lyfter upp en kvinna i en balettföreställning.
I en stad framför en tunnelbana, en man skateboards ner för en trappa som två äldre damer sitter på en bänk titta på honom.
En liten flicka som leker på stranden och bygger ett sandslott.
En liten flicka i gul t-shirt sitter på en sandstrand och leker med sin gröna spade.
En liten flicka glider nerför en tunnel och ler.
En dam som står på trottoaren med bilder på väggen.
Vissa killar spelar basket på en plan.
En man i blå hatt skulpterar en bit is.
Två vackra gröna blomkrukor som sitter utomhus.
En liten pojke går runt med en vit t-shirt och svarta shorts utanför.
Två män dricker öl i en bar.
Två män visas dricka öl medan de sitter i fällbara stolar.
Två berusade vänner dricker en drink till med arga ansikten.
En man i halmhatt och en annan man i randig skjorta som både dricker av koppar och gör roliga ansikten.
Två män gör lustiga ansikten medan de dricker alkohol.
Tre unga flickor går hand i hand i en skara människor.
En man på en motorcykel rider förbi elstolpar och gamla demonterade bilar
En man tar tag i en frisbee medan en annan försöker få den från honom i luften.
En brandman i uniform med mustasch och bock vid sin brandbil.
En samling kvinnor klädda i vitt och rosa på en offentlig torg höja sina armar.
En hejarklackstrupp som uppträder för en publik på ett sportevenemang.
Två personer, den ena rider en vit häst och den andra rider en brun häst.
Folket rider på hästar.
Två personer rider hästar i en tävling med andra människor på hästar i bakgrunden.
En man håller upp en utländsk tidning och tittar på kameran.
En äldre man arbetar på ett fiskenät.
En man som förbereder sitt nät för fiske.
En professionellt klädd man sitter i tunnelbanan och tittar på sin mobiltelefon.
En man som bär mask spelar musik vid sidan av en väg.
En smet gör sig redo att slå bollen kommer mot honom.
En flicka går ner för en gul rutschkana i en pool.
En man målar bokstäver med hjälp av en stencil på en rund stand-up skylt som ligger i sidled.
Mannen som sitter på marken med sitt barn och en barnvagn
En person flyger genom luften på en cykel efter att ha lämnat ett jordhopp.
Det är två personer som deltar i en hästryggsmatch.
Ett band spelar på vad som ser ut som en trottoar snarare än en scen.
En kvinna häller upp drinkar vid ett evenemang.
En äldre man med långt grått skägg sitter på en platt säng.
En man utan skjorta jobbar på ett transportband.
En cykelförare är luftburen från ett hopp medan en annan unge på en cykel tittar på.
Mannen i den blå skjortan jobbar på ljuset.
Flera människor går vid en mänsklig staty, som är målad i olika nyanser av guld.
Två byggnadsarbetare svetsar en metallstruktur.
Unga barn som spelar fotboll på ett frodigt, grönt fält.
Barn som spelar fotboll en solig dag.
En kvinna i grå och blå skjorta ler när hon packar upp och skär i en calzone.
Det finns tre damer klänning i blått stå jublar.
En man och en kvinna som sitter på ett bord på en restaurang och äter middag
En liten pojke som simmar i en pool med mask på.
En svart man i grå tröja och jeans spelar på en gitarr.
En sportkvinna i röd, vit och blå skjorta slutar med en swing.
En ung man i vit hatt spelar golf med en äldre man som bär en blå långärmad skjorta och khakis.
Det är tre personer som plockar grödor från ett fält.
En kvinna, klädd i klänning, sitter ner och spelar ett musikinstrument och sjunger in i en mikrofon.
Tre hanar utför akrobatiska manövrar på en strand medan åskådare tittar på och tar bilder.
En baseballspelare i grå uniform har precis svängt sitt baseballträ på hemmaplan på ett baseballfält.
En lång kö väntar ivrigt på att komma in i ett stängt tält.
Två män tävlar, och mannen framför tittar bakom på den andra ryttaren.
Människan gräver ett blankt föremål ur sanden medan andra tittar.
Två män, en klädd i vita snabels och den andra med röd boxning.
Ett barn sover på en sten mitt i en ånga.
En kvinna i grön skjorta läser en Dr. Seuss bok för tre barn.
Tre män undersöker kläder i en klädaffär.
En cowboy tippar sin hatt med två andra rodeo cowboys, en i en rosa skjorta, en annan i en vit skjorta, båda hästrygg, i aktion, mitt i en rodeo arena.
En asiatisk kvinna vinkar och lutar sig ur en vagn.
En paus i ett tal i Baseball Hall of Fame orsakat av, vad som verkar vara, ett känslomässigt ögonblick.
En gatuarbetare som kör en maskin för att jämna ut den våta betongen.
En kvinna i ett tredje världsland som använder en såg för att skära igenom en stålstång.
Två polospelare rider hästar spelar polo.
En liten hund med ett rött band på huvudet går genom gräset.
En polospelare vaggar en boll medan han rider en häst.
En skallig man i vita solglasögon och en grön skjorta rider en komiskt liten gul cykel.
En man som parasailerar på hårt vatten.
Två killar med blå västar som sitter i uppblåsbara båtar som heter Krossare som är på öppet hav.
En vattenskidåkare vinkar glatt mot kameran.
En rock and roll konsert följer när en gitarrist stjäl rampljuset.
En asiatisk kvinna med ett rött paraply går genom en fullsatt marknadsplats.
Tre män arbetar klädda i orange och gröna uniformer sitter under ett träd för en välförtjänt paus.
En man i vit skjorta doppar en basketboll när en liten publik tittar på.
Denna grupp ungdomar sitter på golvet.
En publik ser två kvinnor cykla nerför gatan.
Cyklister är fokuserade rakt fram när de rider längs en gata med åskådare tittar bakifrån barrikader.
Cyklister tävlar i ett maraton med åskådare tittar.
En fokuserad man bär svart leder flocken i detta cykellopp.
Kustbevakningen är alltid redo att rädda liv i det blå vattnet.
En ung kvinna i blå uniform hjälper en annan ung kvinna i en blå tröja med ett vitt band runt armen.
Två män står och samtalar framför ett flygplan från British Airways.
En kvinna som bär röda leggings och en vit skjorta hänger upp och ner från en metallstruktur.
En man som bär vit skjorta åker skateboard nerför en väg.
Närbild av en cyklist klädd i gult och ridande framför en folkmassa som sitter bakom en röd skylt.
Två cykelcyklister som cyklar utomhus på ett spår.
En kvinna i kostym står på ett podi medan hon talar.
En kvinna kastar champagne på en grupp människor.
Många människor cyklar i hjälmar när fansen tittar och hejar på dem.
En grupp cyklister rider längs tävlingsrutten medan publiken tittar på.
En fotbollsmatch pågår mellan det röda och gröna laget, och det blå laget.
Mannen i rött driver nerför vattenfallet.
En häst och jockey mitt i en hästkapplöpning.
Människor som rider i en Cywedon i cykeldräkter och professionella hjälmar.
Unga kvinnor njuter av utsikten från bron vid lokala festivalen.
Herrarna är på båtdäcket och kopplar av.
En man i blå hatt och orange skjorta lagar en vägs sidospår.
Två barn och en man på en sten.
Lastbilar som omger arbetare mitt på en gata.
En man som ställer in ett skott i snooker.
En kvinna i orange klänning rider på marknaden.
En hockeyspelare i en blå skjorta gör mål mot ett lag i vita skjortor.
Sex hockeyspelare, tre vita och tre blå, skridskor runt det vita lagets mål.
En ung man svävar genom luften på en surfbräda.
Baseball matchen spelas på en cool halv molnig natt.
En man som bär en olympisk fackla med en tegelbyggnad i bakgrunden.
Två män, båda i röda skjortor, en i luften medan de spelar basket.
Två barn som leker på ett metallglas.
En grupp Storbritanniens cyklister försöker trampa sig in i segern.
En grupp simmare hoppar in i en pool.
Två tjejer tävlar och en bär blått är på golvet medan den som bär vitt är ovanpå henne.
En man på en motorcykel som hoppar över en grushög.
En skateboardåkare som bär röd skjorta och knäskydd åker skridskor på en brant ramp.
En dam med gul blus och glasögon vid ett skrivbord med en bärbar dator.
En man i röd skjorta och jeans dansar med en kvinna i en blå och vit klänning på gatan.
Två cyklister tävlar till mållinjen.
Två kampsporter tävlar mot varandra på mattan medan i bakgrunden folk spela in detta och ta bilder.
En ung dam gör sig redo att sjunga in i en mikrofon.
Tre killar i blått och guld njuter av en match.
En grupp cyklister åker ut genom grindarna i en cykeltävling i London 2012.
Fem män i röda skjortor, i en rad, på en basketplan, fyra med händerna på sina hjärtan, och samma fyra tittar uppåt.
En basketspelare från USA dunkar bollen!
Ett lacrosse spel har två spelare i blått och orange spela för ett mål.
En ung blomsterflicka och ringbärare väntar på att få gå nerför gången.
En ung asiatisk kvinna spelar på sin mobiltelefon med sin rygg till sin familj och måltid.
Stolar har placerats framför en byggnad.
Den ekland atletisk spelare försöker vända en dubbelspel som Orioles bas löpare försöker bryta upp det.
En upphängd, uniformerad officer och hans hund går på en strand.
Noggrann hårvård produktapplicering med handske arbetare.
Ett litet barn står på en kulle ovanför en liten fattig by
Tre bicyklister tävlar nerför en livlig gata i regnet, med en röd BMW och en motorcykel som närmar sig bakifrån.
En asiatisk kock tittar på en annan kock på ett galler i ett kommersiellt kök.
I ett område med 2 arméplan, 2 män, en i uniform och en i tunga kläder, träna en svart och brun hund.
Några fotbollsspelare tittar uppmärksamt på bollen och målvakten.
En man i en röd och svart livväst kajaker nerför en fors.
Person med blå skjorta och svart hjälm i kajak i turbulent vatten.
Två kvinnor och en ung man som gräver upp jord och lägger den i en skottkärra.
En afroamerikansk man i marinblått och rött skjuter en basketboll.
En modern sportbågskytt drar tillbaka en pil och siktar.
Fem pojkar i blå skjortor som ritar vid ett bord.
Två Argentina basketspelare, en otroligt glad, och den andra lite frustrerad, med sin tränare klappar för en av spelarna och en kvinnlig chef går från domstolen leende.
En skara olika människor som går genom en marknadsplats.
En man som bär uniform och röda glasögon håller i ett gevär.
En man som lyfter en stor vikt och skriker.
Kvinnlig tennisspelare i gröna shorts och röd skjorta som serverar på en gräsbana på 126 kilometer per timme.
En svettig trummis slår på trummorna.
Trött väg cyklist trycker mot mållinjen som hejas på.
Kvinna poserar i sin monter under London 2012 Olympics
Två patriotiska kvinnor i ryggen av en klassisk cabriolet rida längs i en liten parad.
Folk samlas för Delwood Grannskapets årliga 4:e juli firande.
En hund med vit päls rör sig genom djupt grumligt vatten.
En jockey, ovanpå sin häst, är i mitten av hoppet i en ridtävling.
LeBron James passerar en basket medan bär en USA Jersey medan 4 motståndare står i närheten.
En äldre man sitter på klipporna och ser på när den yngre mannen undersöker vad som finns i vattnet.
Tre män, en klädd i hatt och två som inte är det, knäböjer på marken och gräver i smutsen kring en cementplattform.
En grupp om tre infödda kvinnor vilar i skuggan medan deras barn tittar ut genom en dörröppning.
En man som bär samma färger som cykeln rider nerför gatan.
Två kvinnliga volleybolllag tävlar i ett volleybollspel med åskådare i bakgrunden.
Två lag av kvinnor, en bär blått och rött, den andra bär rött och vitt, spelar volleyboll.
Två tjejlag spelar volleyboll.
Kvinnors volleyboll på OS är mycket intensiv.
Den här mannen har precis avfyrat sitt vapen.
Två personer klädda i fäktningsredskap är svärdslagsmål.
En fäktningsmatch mellan Ryssland och Italien.
Två personer i vita kläder har en fäktningsmatch.
Två unga pojkar leker i sanden nära havet.
En kvinna som bär förkläde och plasthandskar lyfter locket av en bakad vara.
Janitor städar bort dykbrädan med kvast på natten.
En grupp cykelcyklister rider i ett idrottsevenemang.
Flera män i olika färger har en cykel rally.
Två bilar runt ett varv i en professionell tävling.
Tre färgstarka bilar tävlar runt ett spår.
Två staketare, en korean och en amerikan, i en epie bout.
Män i svart och blå springa i bakgrunden som soldat gör push ups i förgrunden.
En man på en surfbräda surfar, medan en stor våg kraschar.
En ung flicka vinkar till kameran medan hon rider på ett ferrihjul.
En kvinna i röd tröja spelar basket.
Brottaren hade övertaget över sin kanadensiska motståndare.
En barfota kvinna, klädd i färgglada kläder, står framför trädet.
En basketspelare bär en vit jersey försöker passera basketen i gränser medan det andra laget blockerar honom.
En person kör en röd och svart racerbil.
En skallig man i en blå skjorta målar graffiti på en vägg
En liten flicka som bär en vit tröja, som sitter framför en färgglad tårta, skrattar med blicken uppåt.
Två kvinnor deltog i en kampsport match innan en publik.
En kampsport turnering i sessionen medan det finns domare i sidlinjen hålla vakt.
En idrottsman springer över tävlingsbanorna på en bana.
Två män hoppar över hinder på en röd bana medan andra tittar och fotograferar dem.
Runners springer längs en bana under ett lopp.
En filmbesättning dokumenterar en kvinnlig idrottsman som kastar spjut.
En målvakt dykning för en fotboll på en fotbollsplan medan kicker klockor.
Två män poserar på ett stenigt område framför ett snöigt berg.
Sex män tävlar under OS i London 2012.
En kvinnlig idrottare använder en kasta anordning för en sport.
Idrottsmän som springer i ett lopp.
En löpare i gröna skor tar ledningen i ett lopp mot en löpare i röda shorts.
Fem unga dam gör sig redo att köra 100m streck
Fyra personer sitter på en sten ute i en vattensamling.
En man i svart hatt som spelar dragspel.
En man rider en häst på en rodeoarena.
En cowboy rotar en kalv i en rodeo.
Två vita hanar spelar squash eller något med en liten boll och en vardera har en paddel.
En man sträcker sig över en annan medan han spelar en sport utanför.
Två kvinnor sitter bredvid varandra, den ena håller ett barn och den andra håller en liten hund.
LeBron James, som spelar för Team USA, försöker lägga sig under korgen.
På en mulen dag, två unga flickor, skratta och leka längs den våta sanden på en strand.
En flicka i VolleyBall-utmaningen, vid OS i London 2012.
Tre flickor är ute i ett sandigt område och spelar volleyboll medan en sittande kvinna i bakgrunden fotograferar dem.
En kanna i röd uniform visas efter att ha kastat baseball.
Två små flickor på en stenväg som håller uppstoppade djur.
En man parasailerar med berg i bakgrunden.
Åskådarna ber att cowboyen inte ramlar av tjuren i rodeon.
Ett barn hoppar över havsvågor vid en strand.
Spelare i ljusgrå uniform når huvudet först för baseballplatta medan catcher i gul topp når armen för att märka honom.
En grupp arkeologer undersöker en utgrävningsplats.
En man med en nummer ett på sin smutscykel åker runt banan.
Detta är en grupp kvinnor som spelar volleyboll i sport bikinis.
Fyra kvinnor i baddräkter som spelar volleyboll på en strand med kameramän som spelar in i bakgrunden.
Fyra kvinnliga idrottare spelar beach volleyboll vid OS i London 2012.
En surfare rider sin surfbräda i början av en våg.
Två män som sjunger i en mörk klubb.
En rallybil bär ner på kameran medan sparka upp en plym av damm.
En kvinnlig idrottsman med nummer 43 på sin kalv springer.
En kvinnlig löpare med solglasögon och grönt med vita sportkläder springer.
En grupp lag tävlar i skogshuggarsporter i British Columbia.
En ung flicka med gunga i ansiktet sitter på ett handfat medan hon gör ansikten i spegeln.
Två kvinnor spelar volleyboll på stranden.
En volleybollspelare som bär en blå bikini förbereder sig för att spetsa bollen.
En ung man förbereder sig noga för att ta en pool shot
Det är två personer som bär solglasögon och hjälmar som står bakom en stor pistol.
Vid ett bord tillsammans med sina kollegor fyller en kvinna i en amerikansk arméuniform i ett diagram.
En flammande rödhårig medelålders kvinna med blek hud står framför en tegelvägg.
Någon, bär en flagga som en mantel, bär 6 öl.
Ett barn mitt på en innergård framför några trappor flyger sin drake.
En vit hund hoppar upp vid en vattenstråle.
En idrottsman rusar nerför en landningsbana som förberedelse för att slunga ett spjut i spår och fält.
En flicka med en enorm hink med blommor.
Det finns en afroamerikansk man som spelar saxofon i en utomhusmiljö.
En man är snål på att gå ombord på stranden.
En man flolics i den gyllene surfing längs en strand vid solnedgången.
En person går i havsvågorna.
En kvinna från Frankrike förbereder sig för att skjuta sin pilbåge med en kvinna från USA bakom sig.
Mannen i orange släppte precis sin pil.
Ett litet barn som håller i en Rawlings-fotboll mitt på ett gräsfält.
En person med röd jacka och längdskidor går uppför ett berg.
Tre barn tittar på groddjur i ett akvarium medan de fotograferar och äter isglass.
Den bas löpare försöker att göra det säkert till väskan.
En ung person färglägger och ritar på trottoaren med rosa krita.
En gentlemän ger en presentation via powerpoint.
Alla människor i parken försöker göra sig bekväma att njuta av programmet som för dem.
En graciös basketspelare står vid den tvåpunktslinjen när hon kastar bollen.
Två killar stannar för att ta en bild medan de håller en flagga.
Mannen hoppar över det andra laget för att spetsa bollen.
En man i grönt ställer in bollen under ett volleybollspel.
Mannen siktar in sig på sitt mål.
En flygman kramar en ung flicka på startbanan.
Två idrottslag tävlar mot varandra.
En man i svart uniform, täckt av lera, drar på sig den lila uniformen av en annan rugbyspelare.
En baseballspelare svänger sitt slagträ för att slå en baseball.
Det finns en kvinna i en blå klänning på den här bilden som verkar resa och väntar på att en tunnelbana ska anlända.
En lacrosse spelare tumlar i mitten av spelet medan andra närmar sig.
En man i jeans och en mörk t-shirt arbetar på ett tåg med en oljekanna.
Racer rider en motorcykel med racerbanan i bakgrunden.
En svart man i blå skjorta spelar en trumma med händerna.
Ung pojke som sitter på en röd sadel på en häst.
Tre kvinnor i rött i det ryska basketlaget jagar basketbollen.
Tre män knuffar vatten från ett baseballfält.
Två personer tävlar i ett cykellopp passerar på vägen.
En grupp reser på baksidan av kameler.
En volleybollspelares solglasögon visar återspeglingen av volleybollen som är framför hennes ansikte.
En guldmedaljör firar sin seger bredvid sin lagkamrat med kameror som omger honom.
Svart och vitt foto av en flicka med korta shorts som springer i regnet med en hoodie på.
En flicka, klädd i en klocka, lagar håret på en annan flicka.
Flera personer arbetar tillsammans i ett skogsområde.
Två kvinnor som spelar basket.
Två byggnadsarbetare lutar sig mot vakträcket på en byggarbetsplats.
Pojke i en flytring i en inomhuspool som tittar på kameran.
Två hanar och en hona sitter vid ett bord på en bar och två dricker öl.
En kvinna som serverar tennisboll.
Flera arbetare klättrar ner för en svagt upplyst tunnelbanetunnel.
En vit kille med solglasögon sjunger med mikrofon.
Två män; en med röd skjorta och fast röd boll, och den andra med en svart skjorta och en lila randig boll, redo att ta en pool skott på ett biljardbord.
En man som bär grå spelar pool i en bar.
En dam med långt brunt hår bär en solbränd tröja och sitter på en soffa med en man.
Mor som håller ett nyfött barn mellan sina morföräldrar medan hon sitter på en soffa.
Stevie Wonder uppträder på scen på en av sina många underbara konserter.
Två unga flickor klappar en liten häst.
En person skär grönsaker på en skärbräda i ett kök.
Motståndsspelare utmanar varandra i ett spel av ultimata frisbee.
En man i gula shorts hoppar i luften för att fånga en frisbee.
Han driver ut sitt hjärta för sitt livs kärlek.
Två män, en med glasögon, simmar bredvid varandra.
Två vita kvinnor som spelar tennis framför en stor publik.
Två bikers, en i svart och den andra med en röd skjorta rida nerför en gata.
Två bicyklister i spandex och hjälmar i ett lopp som trampar uppåt.
En cykeltävling, med cykelförare klädda i flerfärgade uniformer, med en man som spelar in den.
Ett par med slutna ögon dansar när folk ser på.
En olympisk cyklist med nummer 9 från Espania som rider nerför en grusväg.
En manlig badmintonspelare som sträcker sig mot skytteln vid ett OS-evenemang.
En afrikansk amerikansk sångare uppträder på scenen med piano och flera mikrofoner i bakgrunden.
En BMX ryttare i mitten av ett hopp som publiken nedan klockor.
Två kvinnor i långa, ull kjolar är omgivna av getter utanför på en gård.
En man sitter som en man bakom honom tvättar en buss.
Två kvinnor med huvudbonad som pratar i förgrunden med två män i en annan typ av huvudbonad i bakgrunden.
Flera personer med huvudsjalar på en fullsatt marknad.
Stor brun hund som leker med en vit fotboll i gräset.
Två personer fäktas vid OS i London 2012.
En olympisk idrottsman navigerar en slalombana i en kajak och manövrerar försiktigt runt två randiga stolpar.
Olympics kör händelse skjuta från långt borta för att visa den massiva publiken.
Två män med grått skägg delar ett skratt samtidigt som de njuter av det fina vädret.
Världens första och enda skateboardentusiast i Mellanöstern.
En man i en hockeyuniform täckt av annonser som leder en puck ner i rinken.
En flicka som håller upp benet vid sin sida.
En ung kvinna gör en akrobatisk rörelse på ena handen, i en tom pool.
En man kör en smutscykel med nummer 3 på.
Ett litet barn sitter på en matta och leker med ett pusselspel i trä.
En levande spårare vandrar genom en naturskön stig.
En vandrare joggar nerför en stenig väg medan blå himmel och berg korsar horisonten.
En kvinna på en scen möter en fullsatt publik.
En ensam person surfar på en medelstor våg.
En man i en orange kajak paddlar genom stänkande vatten.
Människor i blå uniformer står på gatan när observatörer tittar på från trottoaren.
En man som förbereder sig för att slåss i en basebollmatch.
En närbild av en gitarrist på knä med resten av bandet bakom sig.
En kvinna på en grå och vit häst hoppar över ett hinder.
En man i orange jersey och en kvinna i brunt spelar ett brädspel.
Foursome spelar ett bräde eller kortspel som sitter vid ett bord.
En kvinna och en man öppnar en mixerlåda.
En kvinna laddar diskmaskinen på kvällen efter middagen.
En äldre man i grå tröja och blå byxor formar något i en smedja på ett städ.
Kåken ute på natten går till sin destination.
Flera ungdomar, däribland en ung kvinna i grön och rosa klänning, sjunger och dansar.
Tre tjejer utför en rutin på scenen.
Två unga män utför en modern dansrutin.
Två lag hockeyspelare spelar ett spel.
En man med grått hår sitter vid ett bord.
En man försöker hålla balansen medan han surfar
Tonåringar från olika gymnasier tävlar i en tävling på ett välskött fält.
En grupp idrottare som springer i ett lopp.
En person på en surfbräda med en paddel i en sjö medan två andra människor följer tätt bakom i en båt.
Ett barn i väst och hatt poserar för en bild.
Flickan i rött tar sin tur i Monopol spelet.
En man i grön och vit skjorta och khakis skateboard nära solnedgången.
Den unga pojken i röd och blå dräkt är redo i luften.
Mörkhyade infödda män spelar schack medan de sitter på marken.
Två gröna skjortor fotbollsspelare försöker säkra fotbollen från en spelare klädd i vitt.
Två fotbollsspelare jagar bollen i packade stadion i en tävling mellan USA och Kanada.
En kvinna i rosa skjorta och gul hjälm paddlar runt i en rosa kajak.
En liten flicka och hennes uppstoppade apa satt på en åktur ovanför nöjesfältet.
Tre personer rider motocross cyklar längs en grusväg.
Smutsbiker på en professionell ridbana nära en flygplats, som består av smuts.
Väl ovanför bergens timmerlinje tycks denna unga kvinna vara säkert utrustad för att skala den rena bergväggen.
En bergsklättrare beundrar den vackra scenen i en snötäckt bergstopp.
Bergsklättraren står otryggt på ytan av en stor sten och justerar sin utrustning.
En man uppträder på gatan och spelar två instrument samtidigt.
En surfare gräver sin bräda djupt i vattnet för att skära vågen han rider på.
Ett par tar i utsikten vid vattnet vid skymningen.
Två lag tävlar mot varandra på ett fält i en fotbollsmatch.
En baseball kanna följer genom hans genom.
En man med hjälm på en mountainbike kommer nerför en brant, stenig stig.
En vit kille i svart cykelutrustning rider genom skogen.
Tre personer står utanför ett snabbmatsställe med sina drinkar.
En kvinna sjunger medan en man spelar bongo.
Vacker liten flicka som håller upp sin hatt med ett finger är att få sin bild tagen ut på ett vackert fält.
En kvinna som njuter av en primitiv fläkts vind.
Flickan klädd i rosa bugar sig på ett knä.
En asiatisk kvinna utövar kampsport i en rosa uniform.
Ett litet barn som bär ångkokta glasögon lutar sig mot en grön flytande anordning medan det vilar i vatten.
Två personer tävlar på en BMX-bana.
Fyra paddlare som bär orangea och vita tröjor ro rasande när den sittande publiken tittar på loppet.
En flicka är på trottoaren och tittar på en vit skåpbil på gatan.
En kvinna med en hjärttatuering på sin kalv cyklar förbi ett majsfält.
1 man som cyklar genom landet.
En ung kvinna med bruna byxor rör vid sin sko.
En performancekonstnär upp och nerhängd från röda band.
En grupp människor tittar på ett band som spelar musik medan en dam försöker ta en bild av dem.
En kvinna i ett cykellopp bevakas av en publik.
Bil nummer 14 har kastat upp mycket smuts bakom den.
Det finns ett litet barn, bär en gul flytväst, bär en flytapparat, på stranden.
Tre amputerade i rullstol tävlar tävlingsmässigt på ett spår.
Det är två löpare som just fått köra ett lopp.
Tre löpare är i färd med att korsa mållinjen under ett olympiskt sportevenemang.
En person skalar klippan medan en annan fokuserar på utrustning.
En man som ser mycket trött ut på sidan av en klippa redo att klättra upp till toppen.
En manlig idrottsman i rött och gult dyker mot en badmintonfågel.
En tennisspelare tävlar i OS i London 2012 och hoppar från marken medan han svingar racketen.
En badmintonspelare från Kina är utspritt på Badminton Court med sitt racket i närheten.
Två kvinnor och två pojkar klädda i rosa ställning utanför en butik som säljer färgstarka kläder.
Två små barn går genom högt gräs i skogen.
En matador retar en skadad tjur med sin röda mantel i en turnering.
En man som sjunger och spelar trummor med sin reservgrupp.
Ett team av racerförare i en Ford emblazoned med Mayores förhandlar en sväng på en grusväg.
En racerbil som gör en snabb sväng i ett skogsområde.
En man hoppar med bollen i handen under en plocka upp basketmatch.
En man går för en rebound i en utomhusmatch basket.
En man som har tagit av sig skorna för att knäböja på en matta.
En man spelar ett instrument som omger mina andra män.
En man spelar en handtrumma på sin sista med andra människor i ett band.
En fotbollsspelare hoppar över försvararen.
Två löpare, en svart och en vit, är på banan löper mycket nära i konkurrensen.
En ung dam som sitter på en klippa mitt i en sjö.
En man i utsmyckade stamkläder sjunger mot en fjädrande orange bakgrund.
En pojke njuter av solen, medan människorna i ryggen njuter av havet.
En svart man i blå skjorta håller sitt barn i en blå wrap.
Unge man som åker skridskor medan folk tittar på, i en nöjespark.
En liten flicka i en barnstol har mat över hela ansiktet och fingret i munnen.
En ung person som gör ett högt flygande cykel trick med sina armar ut.
Quarterback Tim Tebow kastar en passning som hans team vakter mot motståndarlaget.
Ung flicka som går över sanden i en blå klänning bär sina skor
En kvinna i en kogirlhatt knäböjer på en hästs sadel medan hon håller handen över sitt hjärta.
Tre personer använder ömsesidiga bankomater från Washington.
En man i blått och en kvinna i vitt dansar med ett annat par som dansar i bakgrunden.
En man fiskar på en bro.
Fem män sitter på ett picknickbord med en skog i bakgrunden.
Människan surfar på en våg i havet
En av medlemmarna i KISS spelar en vit elgitarr framför en svart bakgrund.
En flicka är klädd i en vild outfit dans.
En schäferhund som följer en annan schäfer som har en käpp i munnen.
En kvinna går igenom lite material i en bok med en tonåring.
Person i röd dykardräkt upphängd från en helikopter.
Ett barn, i en blå regnrock, cyklar på en svart väg.
En kvinna med rosa uniform står på en volleybollbana.
En person som kör en gokart svänger till vänster.
En röd bil står parkerad bredvid en svart tjur på ett gräsfält.
En cyklist avrundar ett hörn på en våt väg.
En man i en cykel kastar upp händerna i seger när han korsar mållinjen.
Tre unga pojkar leker med däck, med vuxna i närheten.
Folk spelar vattenpolo och bollen är nära målvakten.
En manlig skateboardare utför ett stunt över en cykel rake.
En grupp människor är utanför och spelar basket medan solen går ner i bakgrunden.
Två staket i full växel tränar sparring.
Två personer som deltar i en fäktningsverksamhet bevakas av en tredje person som sitter på läktare.
En man som sjunger på en mikrofon med rosa skjorta.
Två lag, ett i blått och en gång i vitt, tar sig an varandra för att få kontroll över bollen i detta sportspel.
En umpire som gör sig redo att göra ett nära samtal i en baseballmatch.
En musikalisk artist i en svart klänning berömmer sin publik när röda lampor blinkar och hennes band spelar.
Två konstnärer spraymålar en väggmålning på en betongvägg
En grupp unga blonda barn, en som bär gevär, ställer sig framför ett hus.
Två personer kör i en tävling på ett spår.
Idrottsmannen i körfält 5 spelar in en dominant seger på 2012 års paralympics.
En professionell rullstolstävling med en tydlig ledare i körfält 6.
En grupp kvinnor i mycket dekorerade kläder och silver höga klackar går nerför en gata.
Tre unikt klädda kvinnor som dansar i en parad.
En asiatisk kvinna som ringer står över diskbänken och diskar.
En man bär en svart t-shirt medan han spelar basgitarr i en konsert.
En person som går på en stig med en röd skjorta och blå hatt på.
Spännande åskådare i London hejar på väglöparen.
Kvinnlig ballerina gör en pose upp på tårna av fot i ett stort rum med ett rött golv.
En liten flicka som knyter en liten pojkes sko på gatan.
Männen spelar instrument och pekar på publiken.
En klarröd racerbil kör förbi.
Para-Olympians som representerar Sydafrika i spår och fält fira efter en tävling.
En biltävling äger rum på ett spår.
En man sitter i en fällstol i en bilverkstad medan andra tittar på bilar i bakgrunden.
Två män i tröjor tävlar i en bana och fält atletisk händelse.
Två män paddlar kajak i gula kajaker i ett lopp.
En man i blå skjorta tittar på stenar och träd.
En rodeo tjur ryttare och en hjälpare har mer än de kan hantera i en utomhus rodeo show.
Ett par står på däck på en båt och tittar på vattnet.
En man och en kvinna sitter i slutet av en liten brygga längs vattnet.
Man och ett barn i grå pyjamas leker med en modell bil spår.
Det finns två fotbollsspelare, en bär en blå och gul uniform håller bollen, och den andra bär en vit uniform.
Fotbollsspelare mitt i en match.
En kvinna i röd klänning signerar medan en man i kostym spelar saxofon.
En grupp unga män spelar fotboll.
En skidåkare i blå byxor och röda snöglasögon går baklänges nerför sluttningen.
Två lag tävlar på rullstolsbasket medan de sitter i specialstolar.
En man och en liten flicka skakar hand på spelplanen.
Cheerleaders ordna sig in i en mänsklig pyramid.
Man med lång stolpe som har en korg med eld på spetsen utanför framför två elefanter.
Det här är en ung fotbollsspelare i mitten.
En herrbana möter åtta konkurrenter, alla andra löpare bär orange.
Mor och dotter poserar för ett foto efter att ha vunnit ett pris
En man i vit kostym på en scen interagerar med en liten skara människor som vill ha autografer.
Jackie Chan pratar med kvinnor vid ett OS-evenemang.
En grupp på 7 ungdomar på stranden hoppar i luften och kastar sina skor.
En grupp cyklister tävlar i en tävling.
2 män är klädda i gult och bär halsdukar för att dölja sin identitet, en av dem är levitating över toppen av den andra medan människor tittar på i en upptagen utomhus köpcentrum.
Två män som spelar fotboll på ett plan.
En kvinna hämtar några tallrikar mat från bordet.
Någon kör en klargrön smuts cykel genom gräset.
En dirt bike racer rider nummer 63 över en grusväg i skogen.
Sex mogna asiatiska män som ler mot kameran på sina platser.
En surfare i svart våtdräkt rider vågorna med stranden i fjärran.
En kille som rider en gnarly fem fot våg hela vägen till stranden
Två unga damer kramar kärleksfullt varandra med sina ansikten vidrörande, när de ler mot varandra.
En grupp barn som spelar fotboll vägg sina föräldrar titta på.
Två lag spelar fotboll; det gula hjälmlaget har bollen och avancerar.
En man slår till i en basebollmatch.
En baseballkanna har precis kastat bollen i en hel stadion, det finns en massa fans som bär teal.
En asiatisk man på en tegelgata som tar hand om mat på marken.
En man i blå och svart våtdräkt som seglar i ett blått hav.
Tjej i röd skjorta blåser en bubbla
En tonåring hoppar sin cykel över en ramp framför en gräddfärgad lägenhetsbyggnad.
Tre män står på en plattform.
En skara människor på en stadion utsmyckade i vitt, gult och grönt jubel och klappa för laget nedan.
En grupp människor på en stadion tittar på ett idrottsevenemang.
Folk hejar på fotbollslag på en fotbollsmatch på en stadion.
Detta är en idrottsman på en cykel under ett lopp.
Regal häst och vit vagn scen med kvinnliga förare och två blonda små blommor flickor klädd i vitt.
Kunderna tittar på produkter under en utomhusmarknad av frukt och grönsaker.
En man i vit skjorta har en hög spark med höger ben.
En man är tyngdlyftare med en kettlebell i ett gym.
Bild av 2 cyklister, racing tillbaka till back, förmodligen i motor tvär tävling.
En kvinnlig tandläkare med en äldre manlig patient.
En ung flicka svänger på en gunga framför gräs och träd.
En liveföreställning av två konstnärer.
En pojke leker i en pool med en uppblåsbar leksak.
Två män i röda skjortor tävlar på cyklar, medan andra tittar.
Tre unga pojkar som leker hör inget ont, talar inget ont, ser inget ont
En ung flicka som håller ett boogiebord på stranden
En ung pojke sover på en blå och grön randig kudde på natten.
En familj ber till en utsmyckad staty.
En fotbollsspelare försöker springa runt en på kommande angripare från det andra laget.
ATV racer lutar sig in i hörnet för att upprätthålla sin balans
En ATV ryttare, hastigheter runt ett hörn, medan glider och sparkar upp smuts-fortfarande fokuserad på leden framåt.
En manlig surfare på en vit surfbräda rider en våg.
Två motorcykelförare, med full växel, svänger ett trångt hörn på ett spår.
En person i rött och svart läder som kör motorcykel.
En skäggig man, klädd i jeans och en jacka, förbereder sig för att spela ett flöjtinstrument på trottoaren.
Sex man i en stor kanotliknande båt på lugnt vatten.
På en vacker solig dag, denna unge man utför sporten som kallas vattenskidor.
Ett barn i orange utstyrsel står och håller blommor.
En man som håller i en biljardpinne och spelar pool i ett svagt upplyst rum.
En cyklist rider längs vägen tätt följt av en bil.
En cyklist i rött och svart tävlingsredskap med en aerodynamisk hjälm går nerför en väg.
En blond, kvinnlig fotbollsspelare förbereder sig för att sparka fotbollen.
En baseballspelare som bär vit och röd uniform gör sig redo att slåss under en kväll baseballmatch.
En man och en kvinna på ett produktionsstånd.
En skjortlös man som bär ett korshalsband går bort från en brun tegelbyggnad, med en motorsåg i bakgrunden.
En kvinna med blont hår i röd, vit och blå cheerleading outfit håller vit t-shirt för att svimma.
Spelare från en flickas volleybolllag hukar sig på volleybollbanan.
Racern zoomar förbi skogsområdet och lämnar ett moln av damm.
En äldre man med handskar sitter på en fest nära två kvinnor klädda i kvällskläder.
2 män som tvättar däcket på en båt med en slang.
Två personer är på en klippa med utsikt över havet
Två små barn tittar på trottoaren som de står på
En motorcyklist rusar nerför en tävlingsbana, utan några andra ryttare i sikte.
Unga fans räcker upp händerna medan de lyssnar på en kvinnlig underhållare.
En asiatisk kvinna i hatt mäter mat från tunnor med en slev i en mindre metallpanna.
Kvinnor i hatt en göra säljande varor.
En kvinna sitter i ett marknadsstånd med tre stora brickor med produkter framför sig.
BMX racers rider nerför en brant kulle på en kapplöpningsbana.
En defensiv fotbollsspelare från Wisconsin nästan sparkar UTEP quarterback innan han blev av med bollen.
Kvinnor i Roller Derby är mitt i en match.
Två flickor, på i rött och svart, den andra i blått och gult, spela fotboll.
En man i blå keps och jacka ser frustrerad ut.
En kvinna klädd i rosa är i ett läge med ett ben från marken och en arm i luften.
Ett mycket litet barn bredvid en varuautomat
Två cyklister rider längs en gata i ett maraton som förbipasserande klappar för dem.
Cheerleaders bär vit hålla silver och blå pompoms medan de väntar.
Två kvinnor pratar bakom en bar med flaskor och glasögon i bakgrunden.
En orangeskjortad, manlig golfare, har just avslutat en sving framför en stor publik.
En man i orange och blått har just slagit en golfboll, som en grupp i liknande uniformer ser på.
En man som spelar golf med händerna i luften.
Två killar i ljusblå t-shirts och shorts med vit bokstäver och sport ränder verkar vara igång och aktivt engagerade i ett spel.
En kille i tävlingsutrustning får luft när han rider på en gul ATV.
Många hockeyspelare är hopslagna runt målet, målvakten är i en hukig position och en spelare bär en röd och vit jersey verkar fira.
Två baseballspelare försöker fånga en boll i ytterfältet.
Det finns en cykel showdown så många cyklister ras i en asfalterad väg som åskådare titta på.
En man som cyklade under ett lopp med folkmassor som hejade på honom
En asiatisk bordtennisspelare tittar ivrigt på och väntar på sin motståndare tjänar bollen.
En grupp människor sitter utanför och spelar musik.
Två personer sitter på en bänk lutad mot en byggnad med skrift på den.
En grupp fotbollsspelare försöker ta itu med en annan spelare.
En bild av bicyklister i ett lopp med bakgrunden suddig av deras hastighet.
Någon cyklar i ett cykellopp.
En man i svarta byxor och en blå jacka ser en kvinna sitta på ett trägolv i en brun jacka titta på sex TV-apparater i varierande storlekar.
En ung fotbollsspelare tittar på en match med sin tränare.
Tre fotbollsspelare och en domare hukar sig under en match, medan vuxna tittar i gräsmatta stolar från sidlinjen.
Klättraren försöker bestiga den stora klippan
En flicka i röda shorts går nerför en gata, förbi en byggnad med många gröna växter på väggarna.
En blond kvinna på en spelplan håller sin polosticka redo.
Ett barn i en grön skjorta håller fast vid en axel.
En kvinna som bär en röd blus och en kort står och tittar långt fram
En medelålders man med bruten vänsterarm i kostym, som går förbi ett par kvinnor på trottoaren.
En stor grupp människor i röda uniformer spelar i ett band.
Monster lastbil flyger över gräsiga knolls på en solig eftermiddag.
En man som kör en smutscykel tar en sväng på en stor smutstäckt bana.
I en fotbollsmatch, en Panthers spelare faller framåt i en somersault medan greppa fotbollen.
En fotbollsspelare 94 tar itu med en motståndare.
En fotbollsspelare hoppar över fallna spelare för att fortsätta sin körning.
En fotbollsmatch eller en fotbollsmatch
Manliga fotbollsspelare från två lag går på en fotbollsplan med fans i arenan platser tittar på.
Två hundar slåss om en boll som är i en pöl.
Två män i 60-årsåldern spelar schack i parken
En person med röd skjorta, khakibyxor och en hatt klättrar uppför en bergssluttning.
Två fotbollslag, ett lag bär grönt och vitt, medan det andra laget bär svart, rött och vitt.
Flera män spelar fotboll professionellt utomhus
En arbetare blir utskälld av sin chef i en hård föreläsning.
Den här damen tränar sitt höga hopp på sin nya cykel.
Någon i hjälm som hoppar på en cykel över en stor hög med smuts.
En ung flicka i karatetävling.
En BMX smutsryttare blir extremt hög i luften medan han tittar nedåt på sin nedstigning.
En surfare rider en våg på en stor surfbräda.
Några personer väntar på en tunnelbanestation, med en ankommande bil på avstånd.
En man som surfar i havet.
Ett barn med gumminudel tränas av två män som bär gummiclownnäsor.
En äldre man använder en mountainbike på en stig.
En person som cyklar uppför en grushög medan två andra människor är i bakgrunden och tittar.
Ett synkroniserat simlag som utför en rutin på en tävling.
En vit kvinna, som bär en svart och orange klänning, står framför ett musikstånd.
En orkester som uppträder för en publik.
En man på en cykel faller av den och över en kort avsats.
Petronas racerbil och förare kör på en racerbana.
En gitarrist och trummis är mitt uppe i en liveföreställning.
Gamle skallig man med skägg som sitter ner och spelar flöjt.
Två flickor i vita klänningar står på en kullerstensväg bredvid en vagn och två bruna hästar.
En ung man på en cykling hoppar upp för trapporna på sin cykel.
Människan har sandaler som lutar sig mot ett träd, med andra människor i bakgrunden.
En ung man höjer sin skateboard på en skridskor ramp.
Tre barn är alla leenden när de står bakom galler och poserar för kameran.
Två basebollspelare i randiga uniformer kramas.
Två spelare från New York Yankees kramas medan spelarna runt dem hejar.
En baseballspelare som glider för att fånga en markboll.
En baseballspelare glider in i en bas medan en spelare från det andra laget försöker fånga bollen.
En man med glasögon röker en cigarett.
3 spelare i en fotbollsplan spelar, en tillhör ett lag och 2 i ett annat.
Fyra personer lutar sig mot ett stängsel och tittar på en kulle.
Män spelar ett sportspel med två män i vitt ovanpå en man i svart.
Hockeylagen tar center is för att vända sig mot för kontroll av pucken.
En man sitter på en stolpe framför en dörr bredvid en ikon.
En flicka i ping och en pojke i blått går genom en skogsstig.
Tre killar i uniform lär nio barn att gå med spjut.
De här kvinnorna försöker dansa.
En liten flicka i blå klänning som klättrar på lite gammalt trä.
En ung kvinna i en blå vira runt halsduk sitter i ett museum.
En man i röd skjorta strövar bakdelen av sin cykel i luften vid ett träd.
En liten pojke som leker med nån sorts pipa.
En manlig saxofonspelare spänner ut en sång i ljuset av en lokal anläggning.
Folk går runt på en marknad.
En dam i rosa skjorta som springer en solig dag.
En liten flicka sitter på ett gräsfält med en docka vid sin sida.
En man med en svart och vit rutig jacka och vit färg runt ögonen sträcker sig mot kameran.
En man sitter ensam medan han sminkar sig.
Fotot är på en kvinna i polisuniform som rider på en häst.
En del dansare i mycket färgstarka kostymer som gör en föreställning i ett hektiskt område.
En man på skidor utför ett stunt på ett evenemang med många människor i bakgrunden.
En grupp människor i vita skjortor joggar.
En man i brun rock och byxor står på en fullsatt gata med en blå skylt om Gud.
En indiansk pow wow demonstreras för åskådare.
Snabba fingrar flyger på livliga nycklar som tillhör detta sant att låta Yamaha tangentbord.
En kvinna tittar ut i horisonten medan hon står nära vattenstranden.
Två simmare simmar hals till hals i fristil i simbanor.
Tre personer sjunger och spelar instrument på scenen.
En kvinna på en utländsk strand som håller en matbricka.
En person parasailing över en kropp av vatten och skog område.
Folk festar i en hörsal och en tjej håller upp ett paraply.
En ung flicka i vitt bär en baseballhandske förbereder sig för att kasta en grön boll.
En grupp cyklister färdas förbi en fontän i ett storstadsområde.
En man i röd och gul kostym rider sin cykel genom fältet.
En man med gröna kläder bär sin cykel framför en Rouleur-skylt.
Pilot står bredvid cockpit av flygplan med öppen dörr.
En musiker som håller i en gitarr sjunger själfullt med slutna ögon.
En fotbollsspelare försöker göra mål.
Två barn, en äldre pojke och en yngre flicka, går nerför en trottoar med sina vinterrockar.
En målvakt tittar på handlingen under en fotbollsmatch.
Två unga pojkar är i en brottningsmatch, på en matta.
En tonåring som gör trick med sin favoritcykel.
Ett barn med röda kläder och sandaler i sängen på en smutsig pickup lastbil.
En man i vit skjorta spelar tennis.
En professionell tennisspelare återvänder ett skott med en back hand från ingenmansland.
Den här mannen hoppar på en cykel.
En kvinna i rosa rock står i snön bredvid en "telefonkiosk", och ler när hon håller i en liten spade.
Ett barn står nära ett stängsel.
Lilla flicka i rosa baddräkt hoppar genom en sprinkler leksak utanför.
Två Miami Heat basketspelare har ett roligt samtal.
En man som bär en röd och blå skjorta kör en motorcykel som drar en trailer-last av utrustning.
En kille utan skor som försöker komma på sin cykel.
Fem personer i en gränd nära en rickshaw med en katt som sover på den.
En grupp vuxna spelar ett brädspel vid ett bord
Mannen trummor medan han använder sin öronsnäcka för att hålla jämna steg med musiken.
En ung pojke klappar en katt på en höstväg.
Tre kvinnor som spelar volleyboll och två hoppar för att försöka blockera ett skott.
Två fotbollsspelare som slåss om innehavet av fotbollen.
Två hokey spelare går head-to-head som den förtvivlade kommer undan.
Lilla flicka i en grön barnvagn placerad på runden.
En cyklist bär solglasögon och en silver cykelhjälm tävlar i ett lopp.
Man skär trä inuti en byggnad.
En surfare i en blå våtdräkt fångar en våg medan åskådare tittar i förgrunden.
En kvinna som tittar på något i handen.
En olycklig olycka inträffade på en kapplöpningsbana, där en häst snubblade och föll till marken och tog ner jockeyn också.
Vissa äldre människor spelar ett uråldrigt spel.
En grupp på fyra män som utför en mumlande handling på ett randigt golv i ett mörkt rum.
Vattenpolo simmare tävlar om en lös boll.
En modemodell poserar för kameran med en avslöjande topp.
En kvinna som bär påsar går genom vattnet när hennes hund följer efter.
Två personer går med luffare, den ena är en kort kvinna och den andra är mycket längre och klädd som en clown.
Arbetare sorterar fiskelina.
Musiker på en scen med grönt ljus skiner på dem.
Den skäggige mannen i vagnen applåderar till sina fans.
En ung man i blått och en i bourgogne är i en brottningstävling.
En ung flicka i vit utstyrsel och flip-flops håller två burar
Två kvinnor poserar på en scen med en mörk bakgrund, med armarna upplyfta något.
En man med grått hår bär en solbränd skjorta bläddrar i en samlarbutik.
En man på en cykel rider förbi en park, med en grupp människor i bakgrunden.
En grupp människor står och sitter nära en stor flagga medan de bär traditionella kläder.
I hällregnet ler en maratonlöpare stort när han närmar sig grupper av åskådare, när bilen kör fram bakom honom.
Två löpare är nacke och nacke när bilister rider bakom dem.
En man med nummer 5003 löper längs en gata under ett lopp med hus och mosstäckt vägg i bakgrunden.
En man som är extremt cyklande nerför ett spår.
Två tävlingshästar springer längs banan med nummer fyra före nummer fem.
Folk dansar på en fest.
En man i grå skjorta tar ut två pajer ur ugnen.
Folk dansar i ett rum med en brittisk flagga hängande på väggen.
En grupp unga män och kvinnor som håller i drinkar har roligt i en barmiljö.
Ett par dansar i en tävling med rosa kläder.
Fyra män har kul på Jet Ski's.
En dam i rosa klänning poserar för ett foto.
Två män brottas utan skjortor medan en domare eller domare av något slag börjar lägga sig i.
Utmattandet i kvinnans ansikte medan hon fortsätter att cykla i tävlingen.
En stor grupp tävlande cyklister cyklar nerför en väg kantad av träd.
En liten flicka går en hund vid vattnet.
Två personer spelar gitarr, medan en tredjedel fladdrar trummorna.
Ett nygift par gläder sig bland gästerna.
Fyrverkerier går av, lågt till marken, som folk ser på.
En gravid kvinna som sjunger på scenen medan hon håller en flagga bakom sig.
En kvinna med nummer 697 på tröjan springer i maraton.
En man i röd baddräkt dyker ner i havet.
En man är upp och ner på en utomhusgymnastik bar.
En man och kvinnor kysser varandra.
Två artister, en man som spelar gitarr, och en kvinna med en mikrofon som är upphöjd till hennes mun sitter på stolar som uppträder.
Ett nygift par som skär tårtan.
En man klädd i en jeansjacka som tutar en elgitarr.
En farfar leker med sin familj på en lekplats.
En man gör en yogapose med hjälp av ett träd för stöd i ett stenigt område.
En flicka som bär svart rider en jättestor enhjuling på stranden.
En låg våg bildas i havet mot en grå himmel.
En man i blå skjorta springer.
Fyra män arbetar på en pysselplats med sanden och stranden bakom sig.
Åh, mitt huvud, din dumma a-hål titta på vad du gör nästa gång.
En stående skara människor tittar på en musikalisk föreställning på en upplyst scen.
En man står upprätt på en motorcykel.
Två tjejer sitter på en parkbänk en tittar på sin telefon och den andra tittar på.
Ett lag pojkar spelar fotboll.
En man som springer genom ett fält med nummer 41 märkt på sig.
En ung man står på en gata och håller i en ryggsäck.
En ung flicka med glasögon och svart halsband blåser rök framför kameran.
Tre personer ses på en strand under solnedgången, en hoppar.
En medelålders man i beige väst sover på en träbänk.
Det finns rök framför en tjej med glasögon och massor av halsband.
De unga männen spelar en fotbollsmatch medan mannen i vitt håller mannen i blått.
En familj sitter i en hydda.
Toyota Rally bil plöjer genom en djup pöl av lera på loppet banan.
En tjej som spelar basket i ett gym.
En kvinna springer genom ett fält i regnet.
Hunden springer genom gräset och bär en käpp i munnen.
En äldre man spelar tamburin i en konsert, med en trumpet i knät.
Studenterna förbereder sig för sin banddemonstration.
En asiatisk kvinna är i en rispaddy med kartonger.
En byggnadsarbetare på en dyster dag som skyfflar jord.
Det svarta laget är på väg att förlora mästerskapet mot det blå laget.
En kvinna i fisknätsstrumpor tävlar i en roller derby.
Vid en skateboardpark åker en skateboard, en skoter och 2 man spelar in skateboardåkaren underifrån och ovanför honom.
Två klassiska dansare, en man och en kvinna, uppträder på scenen.
Tre äldre män och en kvinna som sitter vid ett uteserveringshus mot stenmuren.
En surfare som bogseras av en båt har nått en våg.
En man med orange skjorta springer på ett fält.
En liten flicka tittar ut genom fönstret i en tunnelbana.
En grupp människor i sina kajaker förbereder sig för att tävla.
Singer på scen försöker få publiken involverad på en konsert.
En basketmatch med spelare i svart uniform på väg att göra mål medan omgiven av spelare i vitt.
Två små barn leker med färgade bollar.
En man i svart väst spelar gitarr och en annan man spelar gitarr bredvid honom.
En man är klädd i replika ninja kläder.
En rödhårig dam med ett blått förkläde tittar ner på några papper.
Spännande tjejer samlas på en volleybollmatch.
En svart gammal kvinna med grått hår håller fast vid en gul blomma.
Två basketspelare hoppar i luften som en är på väg att göra en slam dunk.
Dirt bike racer i luften med en hand på dirt bike och kropp i luft.
En hornspelare fjäskar framför ett performanceband.
En manlig och kvinnlig vandrare kikar ut över bergen.
Skäggig man bär hatt framför en ofokuserad bakgrund.
Två kvinnor och en man sjunger in i en mikrofon.
Ungdom fotboll spel på en solig dag barn ser runt
Tre barn leker med en boll på en bred gräsyta.
En fotbollsspelare kastar bollen när andra fotbollsspelare tittar på.
En fotbollsspelare springer med bollen och bryter en tackling av försvararen på väg till slutzonen.
En kvinna sitter på en pall och spelar gitarr med ett leende i ansiktet.
En mustachioed man med en rutig skjorta och keps spelar en elektrisk gitarr medan han står vid en mikrofon.
Pojke bär blå kakmonsterskjorta som håller upp ett löv från hösten.
Attraktiv ung kvinna tar en stund att stanna upp och lukta på blomman.
En mörkhårig tjejfärg med orange krita på ett rosa skrivbord.
En man sitter ner och han är omgiven av skor.
En person kryper genom en snötunnel.
En grupp barn som spelar vad som ser ut som violiner i en bandklass troligast i en skola.
Två brottare slåss, brottaren i blått har fördelen.
Tre äldre damer har ätit färdigt på en restaurang och lyssnar på någon som pratar.
En grupp människor som står i en restaurang.
En grupp människor i blått och svart band uniformer med ljusgröna eller röda plymer på sina hattar går genom en publik.
Två barn i blått gör sig av med hästar.
Pojken i de blå shortsen bär en hink på stranden.
En man i vit tröja som står över en öppen grill.
En man klipper bort överflödig lax, så att den kommer att passa bekvämt på en grillplanka av trä.
Två kvinnor, en med rött hår, står utanför en affär.
En dam som kör ett relälopp springer barfota genom lite vatten.
En handfull byggnadsarbetare bygger en mur i ett dike.
En katt tittar på rörelsen av en ung flicka som leker med en leksak flygplan.
Nedförsbacke åkare bär vaddering för att skydda sig när de faller.
Flera män i olika åldrar håller fast vid en bil, medan på skateboards.
Runners tävlar genom knädjupt vatten i ett maraton.
Walkers på en betongpromenad under en blå himmel.
En dam som använder sax att klippa.
En stor grupp unga damer klädda i löparshorts på en startlinje för ett lopp.
En grupp långdistanslöpare tävlar i en tävling.
En basketspelare förbereder sig för att göra ett kast medan hans motståndare försvarar.
En tjej springer med en basketboll, medan en annan försöker stjäla bollen från henne.
En skicklig surfare tar tag i toppen av sin bräda medan rider en våg.
En ung leende flicka i en hatt hukade på ett fält
Ett fotbollslag i gula och svarta uniformer utgör för en bild på fältet.
En svart och vit hund som följer efter några fläckiga gäss.
En del bilar och många tält sätts upp vid foten av ett berg.
En ung pojke som går genom vattnet med ett nät med vågor bakom sig.
En brun och vit hund med en rosa frisbee i munnen sätter sig över en mans rygg.
Folk går runt i ett område med blå sittplatser och en stor tv.
En grupp människor sitter på en soffa och kramar varandra.
Ett ungt par som sitter i en svart stol och ler.
En man och kvinnor smuttar drinkar i två läderstolar.
Folk roar sig på en fest.
Kvinnan som håller upp fyra fingrar har den unge mannens uppmärksamhet i den blå skjortan.
En man framför ett gäng bananer i en svart jacka.
En grupp människor simmar i en flod eller i en liten vattensamling.
Ett barn stänker i havet.
Tre flickor med samma rosa klänning står på stranden och tittar på havet.
Lokala barn leker dragkamp framför en folkmassa.
En man i grön skjorta njuter av en måltid och dricker.
En tjej med en blå och rosa baddräkt som hoppar in i en pool.
En ung kvinna sitter på en bänk och pelar räkor över sin tallrik medan pojken som sitter bredvid henne tar en paus från sin måltid.
En grupp militära hjälptrupper sitter och fyller i pappersarbete i ett rum.
Ett leende barn svingar på en gunga.
Ett professionellt basebollspel som inkluderar The Los Angeles Angels of Anaheim.
En kvinna går för att spela bollen i en omgång beachvolleyboll, medan åskådare titta i bakgrunden.
En dam med svart hår grillar räkor.
En arbetare med ansiktet dolt av ånga från en spis.
En man i vit utstyrsel tvättar en kaklad yta.
En förbipasserande genom att kolla upp vad som finns under spisarnas lock på bordet.
En man uppträder med eldstavar inför en folkmassa utanför.
Ett litet barn hänger upp och ner från en vuxens axel.
Människor som deltar i ett evenemang i en park.
En skidåkare med brun jacka gör ett trick i snön.
Två barn i en inhägnad hundsäng med hunden.
En liten pojke i badkaret spottar vatten.
Kvinna och barn njuta av utsikten från te lakeside.
Två killar sitter i ett rum tillsammans.
Ett barn som rider nerför gatan på en skateboard.
En ung pojke med en stor hatt sträcker sig för att fånga en frisbee.
Två män spelar hästskor.
En ung flicka i röda byxor spelar i ett vattenfontänsområde.
En pojke rider en docka passerade två 1950-tals bilar.
En ung man på en skateboard utför ett trick på toppen av en stenlagd kulle.
Två män klär på sig, och en av dem fixar hans slips.
Studenten sitter i ett klassrum som lärare klädd i gröna föreläsningar.
En man i förgrunden som tränar på en viktmaskin och en kvinna i bakgrunden på ett löpband.
En man med vitt hår, en lång trenchcoat och ett paraply går förbi en parkeringsmätare.
En kvinna går nerför gatan och håller i ett paraply.
Flera personer, inklusive en man i en rosa och svart randig skjorta som tar en bild av något utanför kameran, är i en stads park.
En fårhund samlar ihop en fårhjord.
Ett ungt barn har kul med att leka med en boll.
Ett litet barn i röd skjorta står mitt på gatan.
Två män som bär grå tank toppar och khaki shorts står på byggnadsställningar utanför en tegelbyggnad.
En ung pojke leker med en annan pojke på lekplatsen.
En liten pojke i orange tröja och solglasögon spelar på stranden.
En pojke i rutig skjorta svingar en spade på stranden.
En person står på toppen av en stor, rullande sanddyn.
Arbetare lägger linne i färgat vatten.
Denna thailändska boxare tränar en hög benspark som en uppvärmning innan hans kamp.
En manlig militärläkare ger ett litet barn till sin far.
En man pratar med en kvinna i ett gathörn som bär höga toppar med rosa skosnören.
En liten pojke tittar på fotavtryck i snön.
En man med skägg och solglasögon spelar trummor.
En del människor rider en flotte nerför en vitvattensälv.
Två små flickor ligger på mattan bredvid en O gjord av träklossar.
En traktor försöker plocka upp en annan.
En kvinna och en liten flicka leker med en boll i poolen under några vattenfall.
En man plockar kokosnötter från toppen av ett träd.
En muskulös man som sitter på marken och skär frukt på mitten med en machete.
En pojke i röd kostym hoppar in i en pool.
En man i rutig blå skjorta sover i en stol med bilnycklar i knät.
En man med hatt säljer solglasögon utomhus.
En grupp människor som står på allmän väg, två i förgrunden läser tidningar.
En skara människor vid ett judiskt firande.
En överviktig man och kvinna går på en gata förbi en kaffe &amp; Tea butik.
En koflicka rider på en häst medan han jagar en brun tjur.
En kvinna i cowboyhatt på en häst jagar en kalv runt en smutsring.
Hunden simmar i vattnet
En man arbetar på en jordisk struktur med en pickax.
En man som bär vintermössa skapar keramik.
En man i svart hatt och en blå jacka håller i en hammare.
En man som bär orange skjorta arbetar i ett lerhål
En kvinna i en lång brun rock försöker att cell kvast till två män.
Två män har fullt upp med att tillverka saker i sin butik.
En skjortlös man sitter på marken och håller i frukt.
Två svarta hundar leker med orange objekt kör över gräs.
Flera personer träffas för att spela säckpipa och äta lite mat.
En man som handlar på ett varuhus bredvid en massa godis.
En man med hörlurar arbetar på en laptop i ett svagt upplyst utomhusrum.
Kvinnan sitter på kanten av stockar medan lugnt ligger i ett risfält.
En man visar en ung pojke hur man sopar på gatorna i en asiatisk stad.
Två män skriker åt en kvinna på en marknadsplats.
En man i en svart långärmad T-shirt ser fram emot att prova lite mat som har lagts ut på ett soffbord.
Ung blond kvinna sätter sin fot i en vattenfontän
En tygarbetare tittade uppmärksamt på kameran och pekade på honom.
En man i röd hatt som böjer sig över.
Två pojkar med blont hår, klädda i randiga skjortor på en säng.
Flera barn klättrar stora stenar i en park.
Svart hund med krage hoppar upp med en pinne i munnen
En asiatisk gatuhantverkare modeartiklar till salu.
Tre män arbetar för att förtöja en stor båt till kajen.
En Zoo-hanterare ägnar sig åt en aktivitet med en vit tiger.
En pojke som bär mörka kläder ligger på en röd filt vid tältets öppnande.
En liten pojke leker i en sprängleksak.
Tre personer i ett rum med en kvinna i svart skjorta och hals halsduk som håller en drink i handen.
En man i gul skjorta inspekterar smycken i en smyckesaffär.
En man med vit skjorta och blå byxor som lagar en hälsosam måltid med grönsaker.
En pizzakock koncentrerar sig på något.
En kvinna läser en annan kvinnas handflata vid ett blått bord.
En mörkhårig kvinna sätter en etikett på en cigarr.
Två damer gör klart för servering.
En familj poserar med SvampBob Squarepants.
Människor som passerar genom en öppen marknad, medan en äldre kvinna lutar sig framför en kyld bin on=f skaldjur.
En byggnadsarbetare balanserar på en byggnadsställning.
Det finns en man som arbetar på en tårta dekoration med ett litet, tunt verktyg för att hjälpa honom att skapa intrikata former och mönster.
En man med skägg i coveralls på en skaldjursmarknad.
Damen med håret upp i en bulle, i en tank topp och khakis tittar på ett starkt ljus.
En reporter pratar med en kvinna medan åskådare tittar.
En ledare i overall och en blå hatt står utanför en bil i ett lokomotiv.
En fönsterputsare balanserar sig själv medan han torkar fönstret.
En herrar i en bourgogne långärmad skjorta är på ett fruktstånd som säljer vattenmelon.
En mycket glad ung kvinna som lagar ett mellanmål.
En man går igenom sin skrotbok och beundrar minnena från sina resor till Kina.
Två män på en körsbärsplockare sätter upp en skylt med en kvinna.
Tre kvinnor och en man klädd som "naken cowboy" i New York.
En liten pojke i blått som gör cykelhopp.
Ypoung flicka med armar korsade över hennes hjärta bär en bikini inställning i högt gräs framför en kropp av vatten.
Två män rusar hästar under en rodeo.
En man som bär cowboyhatt, rider på en bronco medan en annan man i vit skjorta kommer till hans hjälp.
Damen med kundvagnen är omgiven av leksaker galore och olika barncyklar.
Fyra barn tittar på TV medan de sitter i stolar.
Två män äter mat i en cafeterian.
Fyra unga män som håller i koppar och mat är i en kurragömma.
Två personer går förbi en industribyggnad.
Gatuförsäljare med Nescafe vagnar pratar med varandra i ett hörn med julgranar.
Två damer säljer frukt och producerar på gatan.
En underhållsarbetare på händer och knän som rensar ut dräneringsdiken.
En man vilar sitt huvud på bordet med slutna ögon.
En grupp människor går medan de håller många korgar och mattor.
En skäggig man sitter vid ett bussfönster.
En grupp bilder i ramar arrangeras med färgglada blommor placerade framför dem.
En tjej i vit skjorta och kjol som spelar tennis.
En man dammsuger en matta medan ett litet barn trycker på ett leksaksvakuum bredvid sig.
En ung pojke skjuter ivrigt en basketboll.
En publik tittar på när flera kvinnor drar på ett rep, kanske spelar bogserkrig.
Två barn spelar hockey på en damm.
En kille med gyllene hår pratar med en kille med rött hår på huvudet.
Två kvinnor tar hand om vissa djur.
Dessa två cykelcyklister njuter av en stig längs en flods kant.
En man förbereder en varm dryck.
En man med håriga armar och en klocka häller grädde i en kopp kaffe, gör färg krusningar längs ytan.
Två kajakpaddlare; en paddling och en i vattnet.
Morfar visar hur den stora gula borren fungerar så att pojken vet hur man hanterar den orange leksaks borren.
En ung asiatisk flicka med en vit björnstrumpa.
En lärare och hennes elever är i klassrummet alla bär vinterjackor.
En artist som visar upp sina färdigheter på en show.
En man sitter bredvid en massa material medan han syr.
En gammal man står bredvid ett skruvstäd.
En man i blå skjorta och en ung flicka i lila skjorta i ett torrt, stenigt område.
Lyckligtvis prövar en ung kvinna sin nya repsving.
En man med en färgstark hatt sitter bredvid en mängd olika verktyg.
En man överväger sitt nästa drag när han bygger om sitt utrymme.
En man med lång maroonhatt trummar på en svart metallskål.
En kvinna spelar gitarr för två små barn.
Mannen läser för sin son medan mamma tillbringar tid med det andra barnet i soffan.
En kvinna som bär en rosa Tinker Bell-jacka lutar sig mot ett räcke.
Två pensionärer tittar som en liten pojke flolics och pjäser.
En clown klädd i rött och gult håller något i munnen.
En man i bredbrydd hatt sover mot en pelare.
Två män och en kvinna är i en inspelningsstudio.
En svart hund står ovanpå en brun hund på gräset.
Många människor sitter eller står runt fontänen nära Space Needle.
En tjej i en rutig, grön skjorta som hoppar i luften.
En man klättrar uppför ett berg.
En pojke i flytväst hoppar på något gult, utom ramen.
Fem byggnadsarbetare bygger en grå byggnad.
Två kvinnor äter av flera vita rätter.
En man som bär ryggsäck hoppar från en pier.
En man i gul kort och shorts jonglerar knivar.
En hund hoppar i gräset.
En dam med röd skjorta som håller en kopp smaksatt is.
Kvinnor i kostym står på en scen.
Två unga män arbetar över en grill och lagar och serverar mat på käppar.
De två kvinnorna och pojken sitter.
En man sitter ensam på en soffa i ett timmerrum.
En man i halmhatt målar.
En grupp män på trappor som leder till en stor vattenförekomst.
En brud skrattar när en äldre man talar in i en mikrofon.
Två kvinnor i bikini spelar bordtennis på stranden medan en annan kvinna i en handduk klockor.
En vit hund springer längs stranden
Två brandmän från Aurora har ett samtal framför en butiksfront.
Ett gift etniskt par firar bland kamrater.
En liten pojke i en taupetröja försöker fånga en grön ballong ovanför honom.
Flera barn är runt ett bord med en ljusblå duk.
Flera kvinnor går nerför gatan klädda i rosa och andra blandade människor.
En man och en kvinna står på ett fält.
En man i en folkmassa håller kamerautrustning som om han är på väg att ta en bild.
En äldre kvinna som säljer ris på gatan.
Folk är i ett kök, två av dem sitter vid köksbordet.
En diskjockey blandar musiken när tjejer dansar bakom honom.
En kvinna i en tank topp sitter och stickar vid ett bord, med en flaska av något att dricka bredvid henne.
Två kvinnor drar i en annan kappa.
En kvinna slappnar av i en utomhus spa på omgiven av majestätiska berg och breda öppna dessert fält.
Den här flickan lägger fågeln i snö, och äter den senare.
En person hänger i ett säkerhetsrep när han klättrar ner för en stor klippa.
En kille med ett gult armband som skär i en tårta.
Två män sitter på en flygplats och väntar och skriver i anteckningsböcker.
En flicka som täpper till näsan under vattnet.
En kvinna med grå byxor, blå skjorta och sneakers sitter i en stol och skriver på en pad.
Två unga män spelar trumpet i traditionell mariachiklänning.
Tre personer i blonda peruker och svarta klänningar som sjunger till mikrofoner.
Mannen går med ett litet barn utanför.
En man och en ung pojke som sover i en stol.
En grupp pf personer som är närvarande vid ett firande
En grupp människor cyklar på en gata.
En person i luften som gör en backflip.
En hund hoppar upp på bakbenen med munnen öppen.
En man i blå skjorta skär i träet.
En pojke i svart baddräkt som leker nära vattnet.
En kvinna som pratar på en mobiltelefon inne i ett stort byggnadskomplex.
Mannen i den röda skjortan klättrar upp på sidan av ett berg.
En bror och syster tar en stund att fnittra och ha kul under karateträningen.
Pojke och flicka som övar marskalkskonst på en blå matta.
Två vuxna leker på ett barnpass.
En man har en stor fisk på en båt.
En grupp män gör husreparationer.
En man i svart hatt står bredvid en svart stolpe.
Brandmän sätter eld på oss.
Brass-sektionen i en orkester, mestadels i skolåldern, framför ett stycke.
Tre barn klättrar upp på ett boskapsstängsel.
En man med glasögon och en långärmad grön skjorta beundrar en Komodo drake.
Barnet försöker dricka från två sippiga koppar.
Kvinna i vit skjorta och blå och vita shorts promenader.
En hund springer genom ett fält och jagar en boll.
En ung pojke drar en annan pojke med en fånig hatt i en radioflygvagn.
Barn som simmar under vattnet med en leksak i handen.
En kvinna som knådar deg i köket med bara händerna.
En man häller smet ur en silverskål.
En man tar en bild av något man inte ser till höger.
En kvinna som springer efter ett barn på stranden.
En man klättrar upp för en mycket stor sten.
En ensam båt som sitter i vattnet.
En man i brun t-shirt och blå jeans står framför en chanelbutik och håller en walkie talkie.
En man lagar mat på en grill utanför ett hem.
En äldre man står ensam i kostym och slips utanför en affär.
Tre små pojkar med nät som letar efter insekter att fånga.
Framför finns en kille som sjunger och spelar gitarr och en vit tröjad trummis på baksidan.
En liten flicka springer genom inkommande surfing på en strand.
Asiatiska skolbarn sitter på varandras axlar.
En man i en brunfärgad skjorta skär mat.
En man med glasögon sitter vid ett skrivbord och håller i en telefon och några papper.
En man som vilar i en grunt flod mitt i klipporna.
En fiskare står på några klippor vid havet, upplyst av solen, som är nära horisonten.
Baseballspelare tittar ut i en stadion publik
En turist går nerför gatan, kamera i hand, försöker hitta något värdigt ett foto.
Sju vuxna sitter vid en brandstation och pratar.
En pojke hoppar över en blå slangpipa som en liten flicka klockor.
En liten hund i koppel känner lukten av ett annat djur.
En kvinna i vit skjorta och glasögon målar en vit vägggrön.
En pojke klädd i röda krokodiler som klättrar upp i ett träd.
En flicka som bär orange skjorta håller i stolpar och tittar ner.
Ett rum fullt av folk som äter vid runda bord.
En man med glasögon och en vit klänning skjorta sitter längs sidan andra kvinnor och män på en middag.
En kvinna knäböjer nära vattnet.
En ung pojke står bakom en vävd matta under ett tak av palmfronder.
Man spelar elgitarr live under en konsert.
En kille i blå jeans med svart skjorta har handen i fickan.
En ung flicka knuffar en leksak medan hennes tvillingsyster ser på.
Två män och en kvinna sitter vid ett bord och äter efterrätt.
En hane klipper gräset med en gräsklippare.
Den gula hunden dricker vatten från en flaska.
Tjejen simmar i en sjö under vattnet.
En pojke i en ljusblå t-shirt och röda shorts springer framåt när han svingar ett basebollträ bakom honom.
Folk åker skridskor och går över en frusen yta med Adobe-byggnaden i bakgrunden.
En kille i svart jacka och blå jeans håller ett stort arrangemang av rosor medan du går längs trottoaren.
Två flickor sitter bredvid en flod under ett träd
Någonstans i en varm dessert några människor går med och några på hästar.
En ung pojke står på trottoaren medan en man lyfter upp en väska i bakgrunden.
En liten hund hoppade kastade lite en sjö
Man och ung pojke sjunger tillsammans med mikrofoner.
En man i jeans och en lila skjorta hårt på jobbet bygga en däck.
Isskulpturer får en helt ny innebörd i Alaska.
En man går förbi träd framför stadens skyline.
En hundvalp leker med en tennisboll.
En man i svart skjorta njuter av ett mellanmål medan en kvinna i vit skjorta ser förvirrad ut.
En ung man som sitter och klappar sin hund
Grupp av människor under fana med symbol på den.
En grupp människor förbereder en varmluftsballong för flygning.
En person i en svart jacka mitt på vägen.
En man med rutig skjorta, grädddräkt och tennisskor sitter på en bänk.
En kvinna med glasögon som ska ta en tugga av en stor kaka.
En pojke poserar för ett fotografi på stranden.
Barnet som bär mössa håller i en fiskespö.
En man i idrottskläder inspekterar en svart och röd cykel.
Två män städar utsidan av en byggnad under en blå himmel.
En liten bebis sitter på en säng och ler.
En tjej i en blå gymnast outfit hoppar och gör delar.
En man i fiskeoveraller i vattnet.
En ung, blond flicka står utanför och blåser bubblor.
Ensamma skidåkare går genom snön.
Ett marschband i röda och vita uniformer.
En kvinna klättrar uppför en klippa
En kvinna med hatt som säljer något till en äldre kvinna med vitt hår.
Tre pojkar leker längs en inredningsvägg utanför en byggnad.
En man i blå jeans och en ung pojke i brun skjorta leker i trädgården.
En grävsko gräver ut smuts i skymningen.
En kvinna som drar en vagn med en flicka i den över en frusen sjö
En skäggig man med djurhudsrock och hatt.
En flicka sitter vid ett bord framför en tallrik mat.
En äldre kvinna vänder sig bakåt och skriker.
På liknande sätt spelar barnen fotboll på ett stenigt fält framför en byggnad.
En svart kvinna med hatt på väger frukt och grönsaker.
Flera beskyddare står ute i regnet för att få tilltugg från en gatuförsäljare.
En pojke och en hund står på en brygga och tittar på en annan hund.
En man med glasögon på och en bandanna som täcker hans mun tittar ut genom ett fönster.
En person sitter under ett lila paraply på stranden.
Ett litet barn står framför en spegel och har svårt att ta av sig sin röda jacka.
Flickor i baddräkter, håller i händerna och hoppar ner i vattnet.
En ung pojke i gul skjorta leker med lite utrustning.
En liten flicka med uppblåsbara armband hoppar in i poolen
En svart hund med röd krage har ett föremål i munnen och klättrar upp ur en pool.
En man sitter framför en bankomat medan en annan man använder maskinen.
En man med vit hatt sitter vid ett bord och lyssnar på en man som sjunger och spelar gitarr.
En grupp gamla män samlas runt en bil.
En kvinna klipper ett får på ryggen framför en röd tegelvägg.
En kvinna i tröja rör vid ett får.
En brunhårig kvinna knäböjer medan hon samlar ull på en svart presenning.
Man i röd skjorta klättrar klippa
Kvinnan i blått kastar ett litet barn i en pool.
En man som sitter på en stol bredvid böcker sover.
En man i solbränd jacka och blå jeans sitter och tittar på pappret.
Ett bergslandskap.
En ung flicka i rosa jacka bär en rullande bagageväska
En man i hatt går på en parkeringsplats.
Två personer gör sitt jobb bra och visar upp sig för allmänheten.
Människor gör olika aktiviteter i en park.
En pojke i gul t-shirt leker med en leksak som liknar en dammsugare slang.
En stor publik tittar på något slags spel.
En beagle som går på stranden bredvid några vågor.
En kvinna som bär en rosa tanktopp som håller i en mugg vätska
En kvinna som jobbar på en vinbar och bär ett vitt förkläde.
En kvinna som gör smutsiga handarbeten på trä.
En löpare med en grön sko och en vit sko springer uppåt.
En man i en solbränd jacka sjunger in i en mikrofon.
En pojke slickar en äldre mans ansikte som är täckt av ett blått och gult krämigt ämne.
Man rider cykel på spåret
Två män sitter mot ett stenmonument bland snötäckta toppar.
Det finns två män som cyklar utomhus på den snötäckta landsbygden.
En man på cykeltur högt uppe i bergen.
Mannen på cykeln sitter på en gruskulle.
Fyra personer tittar på något på väggen i ett väntrum.
Två hundar brottas på ett fält.
En vandrare navigerar ett rep och en träbro över en stor torr ravin.
En man tar en tupplur på tåget.
En man i vandringsstövlar, shorts, en blå jacka och en bred brättemössa går genom ett område med tallar.
En ung man som står på en uteplats.
Solstrålar lyser ner på ett grönt tält i skogen.
En man och en kvinna gör en akrobatisk pos i en pool.
En man i hatt målar ett trästaket utanför.
En mässa i Texas med många människor.
En ung blond pojke sitter i slutet av en brygga och håller en fiskespö över vattnet.
Par samlades i en brickbyggnad som gick nerför trapporna.
En kvinna i vitt och en man i svart kostym skär tårta tillsammans.
En far med sin son som gick på gräsmattan.
En man som tar på sig geisha som smink i en spegel med en vit skjorta
En väldigt smutsig ung blond pojke som leker i leran.
Ett lag i gula, röda och blå tröjor sitter bredvid en väg och tittar på en tiger maskot.
En ung flicka med en tutudans i ett stort rum.
En grupp människor som bär ljusblå skjortor och mörkblå byxor som rör sig runt alla tillsammans.
En liten pojke som bär en vit skjorta trycker på en grå kundvagn.
En kvinna med en svart väska som väntar på en orange busshållplats.
En matsal full av människor som äter och en servitör som serverar dem.
Två män försöker driva denna mycket stora uppblåsbara golfboll
Ett barn leker med en leksak i gräset.
En man i röda stammar flyger genom luften med en boogiebräda.
En grupp ungdomar som pratar och skrattar.
Två kvinnor och en man är i en sportig röd cabriolet framför en stor grupp människor på trottoaren.
En kvinna som sover ensam i en säng.
Två rörpassagerare svetsade en söm vid en stor koppling.
Mannen håller ett barn nära en karneval spel.
En man som ler in i kameran samtidigt som han håller en dekorativ platta och en bläckpenna
Ett par kysser högst upp på trappan på en trottoar.
Fyra unga vuxna med två mikrofoner gör dumma ansikten vid kameran.
En hund hoppar ner i vattnet nära en motorbåt.
Två pojkar klättrar upp i en träplattform och hoppar ner i en flod.
Ung flicka som bär en baddräkt med två delar som badar under ett litet vattenfall.
En liten flicka med lockigt hår med öppen mun.
Den här killen, vit skjorta, och blå Shorts tar en sväng någonstans.
En brun hund springer över snö nära lövfria träd.
En man med smutsiga fötter som ligger på ett steg utanför.
En del vandrare korsar en trä- och trådbro över en flod.
Personen går i bergen.
En grupp människor som står på en balkong i en mycket modern miljö.
En pojke i grön skjorta gör en haka uppåt.
Två män i traditionell arabisk klänning står nära en bil våg vid en SUV i öknen.
Människor som sitter inne i en buss och väntar på att nå sin destination.
Simmare hoppar från startblocken in i sina kapplöpningsbanor vid en inomhuspool.
En man som just kom från ett bad.
En kvinna använder en symaskin för att sy på sidan av gatan.
En kvinna med rakat huvud klädd i svart och vitt i en parad
Två barn, en hane och en hona tränar utomhus bergsklättring.
En äldre skäggig man som vilar i en förfallen byggnad.
En kvinna kastar vatten på ett barn i en plastpool på landsbygden.
En hund och en katt slåss på en stol.
Ett barn som leker med en vattenslang medan en kvinna spelar in med en videokamera
En man som sitter ner njuter av sitt kaffe på ett kafé.
En liten pojke klappar en tiger som ligger ner.
En man klättrar uppför ett isigt berg.
Två personer sitter i fjärran på en ovanlig klippformation.
En grupp människor går nerför en trottoar.
En kvinna i en labbrock tittar genom ett mikroskop.
En medelålders, lättklädd man rekvisiterar sina fötter på sitt skrivbord.
En vagn innehåller två män som dras av hästar i regnet.
En vit liten flicka kramar en svart kvinna.
En etnisk gatuförsäljare ler när han visar upp sina grönsaker och röker en cigarett.
En långhårig hund med rosa väst och löpning
En man i blå jeans och en vit t-shirt arbetar på ett fönster med rälsvakter.
En indisk man pratar med barn när de skär en tårta.
Två kvinnor i baseballmössor står mot varandra i en fullsatt hörsal.
Ett barn sjunker ner från vattnet.
Två flickor går bort från kameran under en gångväg.
Sex små barn sitter vid ett skrivbord.
Judiska män och pojkar som sitter och läser Torán.
En möbelaffär har samlat en stor mängd människor.
Ett litet barn i röda och svarta vinterkläder står nära ett stationärt tåg.
Människor som står med tecken som representerar fred i sina händer.
En kvinna visar ett fredstecken medan hon står bredvid ett barn som håller ett ballongdjur medan hon äter mat på McDonalds.
En grupp människor som går vid en sjö.
Byggarbetare står på baksidan av en sopbil.
En äldre kvinna som sitter i ett kafé och har en jacka och läser en bok.
Två vita och bruna hundar mot ett staket.
Två män använder verktyg på det här trädet.
En manlig polis skriver en biljett bredvid en bil.
En säckpipa street artist framför ett skyltfönster.
En man och kvinna som håller träundersökningar och utövar kampsport rör sig framför en folkmassa.
En grupp män sitter ner på marken tillsammans.
En pojke glider ner i en röd skjorta.
Ett asiskt par njuter av sushimiddag
En grupp solbadare ligger på klipporna på handdukar och filtar.
En person går med en vit väska.
En kvinna i en röd blommig klänning med cardigan tar ett foto på en naturstig samtidigt som hon håller ett regnbågsparasoll.
En man och en kvinna gör sallader.
Två män övar kampsport i en trägolvsstudio.
En man i karate poserar på ett trägolv.
Folk står utanför caféet och ska gå in.
De två hundarna springer genom gräset.
En fabriksarbetare tar en paus från sin dag för att posera för kameran.
En pojke i vinterkläder glider ner för en orange rutschkana.
En person bär på en spade som går nerför en snöig gata.
En flicka i gröna glasögon i en pool med tre andra barn.
Den svarta hunden har en leksak i munnen och en person står i närheten.
En man gör en wheelie på en mountainbike.
Tre män, en med skorna av, sover på en bänk i parken.
Fem personer sitter tillsammans i snön.
En kvinnlig gymnast i en svart endräkt och beskådas bakifrån förbereder sig för ett tumlande pass.
En kvinna på golvet täckt av tårta.
En polis som stod på gatan tillsammans med tre poliser på hästryggen.
En kvinna talar på ett podi utomhus.
En äldre man håller en burk bakom ryggen när han promenerar förbi en vacker blomstermarknad.
En man som sätter ihop en trästol.
En grå fågel står majestätiskt på en strand medan vågorna rullar in.
En man i silver regnrock står utanför vid en skottkärra.
En kvinna bakom en rulled vägg skriver
En bergsklättrare övar på en bergsklättringsvägg.
Två manliga byggnadsarbetare arbetar på en gata utanför någons hem
En äldre man sitter utanför en butikslokal tillsammans med en ung pojke med en vagn.
En man i shorts och en Hawaiisk skjorta lutar sig över rälsen på en lotsbåt, med dimma och berg i bakgrunden.